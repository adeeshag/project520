
module updateY_datapath ( clock, reset, executeEnableBit, yInVal1, yInVal2, 
        op_yWriteVal, op_DoneFlag, op_ExDoneFlag, op_CPDoneFlag, op_fpIn1, 
        op_fpIn2, op_fpMode, in_fpOut );
  input [47:0] yInVal1;
  input [47:0] yInVal2;
  output [47:0] op_yWriteVal;
  output [47:0] op_fpIn1;
  output [47:0] op_fpIn2;
  input [47:0] in_fpOut;
  input clock, reset, executeEnableBit;
  output op_DoneFlag, op_ExDoneFlag, op_CPDoneFlag, op_fpMode;
  wire   U17_DATA2_0, U16_DATA2_0, U11_Z_0, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n574, n671, n672, n673, n674;

  SDFF_X1 op_ExDoneFlag_reg ( .D(n55), .SI(1'b0), .SE(n164), .CK(clock), .Q(
        op_ExDoneFlag), .QN(n50) );
  DFF_X1 op_DoneFlag_reg ( .D(n54), .CK(clock), .Q(op_DoneFlag) );
  DFF_X2 temp_yComputedVal_reg_47_ ( .D(n207), .CK(clock), .QN(n2) );
  DFF_X2 temp_yComputedVal_reg_46_ ( .D(n208), .CK(clock), .QN(n3) );
  DFF_X2 temp_yComputedVal_reg_45_ ( .D(n209), .CK(clock), .QN(n4) );
  DFF_X2 temp_yComputedVal_reg_44_ ( .D(n210), .CK(clock), .QN(n5) );
  DFF_X2 temp_yComputedVal_reg_43_ ( .D(n211), .CK(clock), .QN(n6) );
  DFF_X2 temp_yComputedVal_reg_42_ ( .D(n212), .CK(clock), .QN(n7) );
  DFF_X2 temp_yComputedVal_reg_41_ ( .D(n213), .CK(clock), .QN(n8) );
  DFF_X2 temp_yComputedVal_reg_40_ ( .D(n214), .CK(clock), .QN(n9) );
  DFF_X2 temp_yComputedVal_reg_39_ ( .D(n215), .CK(clock), .QN(n10) );
  DFF_X2 temp_yComputedVal_reg_38_ ( .D(n216), .CK(clock), .QN(n11) );
  DFF_X2 temp_yComputedVal_reg_37_ ( .D(n217), .CK(clock), .QN(n12) );
  DFF_X2 temp_yComputedVal_reg_36_ ( .D(n218), .CK(clock), .QN(n13) );
  DFF_X2 temp_yComputedVal_reg_35_ ( .D(n219), .CK(clock), .QN(n14) );
  DFF_X2 temp_yComputedVal_reg_34_ ( .D(n220), .CK(clock), .QN(n15) );
  DFF_X2 temp_yComputedVal_reg_33_ ( .D(n221), .CK(clock), .QN(n16) );
  DFF_X2 temp_yComputedVal_reg_32_ ( .D(n222), .CK(clock), .QN(n17) );
  DFF_X2 temp_yComputedVal_reg_31_ ( .D(n223), .CK(clock), .QN(n18) );
  DFF_X2 temp_yComputedVal_reg_30_ ( .D(n224), .CK(clock), .QN(n19) );
  DFF_X2 temp_yComputedVal_reg_29_ ( .D(n225), .CK(clock), .QN(n20) );
  DFF_X2 temp_yComputedVal_reg_28_ ( .D(n226), .CK(clock), .QN(n21) );
  DFF_X2 temp_yComputedVal_reg_27_ ( .D(n227), .CK(clock), .QN(n22) );
  DFF_X2 temp_yComputedVal_reg_26_ ( .D(n228), .CK(clock), .QN(n23) );
  DFF_X2 temp_yComputedVal_reg_25_ ( .D(n229), .CK(clock), .QN(n24) );
  DFF_X2 temp_yComputedVal_reg_24_ ( .D(n230), .CK(clock), .QN(n25) );
  DFF_X2 temp_yComputedVal_reg_23_ ( .D(n231), .CK(clock), .QN(n26) );
  DFF_X2 temp_yComputedVal_reg_22_ ( .D(n232), .CK(clock), .QN(n27) );
  DFF_X2 temp_yComputedVal_reg_21_ ( .D(n233), .CK(clock), .QN(n28) );
  DFF_X2 temp_yComputedVal_reg_20_ ( .D(n234), .CK(clock), .QN(n29) );
  DFF_X2 temp_yComputedVal_reg_19_ ( .D(n235), .CK(clock), .QN(n30) );
  DFF_X2 temp_yComputedVal_reg_18_ ( .D(n236), .CK(clock), .QN(n31) );
  DFF_X2 temp_yComputedVal_reg_17_ ( .D(n237), .CK(clock), .QN(n32) );
  DFF_X2 temp_yComputedVal_reg_16_ ( .D(n238), .CK(clock), .QN(n33) );
  DFF_X2 temp_yComputedVal_reg_15_ ( .D(n239), .CK(clock), .QN(n34) );
  DFF_X2 temp_yComputedVal_reg_14_ ( .D(n240), .CK(clock), .QN(n35) );
  DFF_X2 temp_yComputedVal_reg_13_ ( .D(n241), .CK(clock), .QN(n36) );
  DFF_X2 temp_yComputedVal_reg_12_ ( .D(n242), .CK(clock), .QN(n37) );
  DFF_X2 temp_yComputedVal_reg_11_ ( .D(n243), .CK(clock), .QN(n38) );
  DFF_X2 temp_yComputedVal_reg_10_ ( .D(n244), .CK(clock), .QN(n39) );
  DFF_X2 temp_yComputedVal_reg_9_ ( .D(n245), .CK(clock), .QN(n40) );
  DFF_X2 temp_yComputedVal_reg_8_ ( .D(n246), .CK(clock), .QN(n41) );
  DFF_X2 temp_yComputedVal_reg_7_ ( .D(n247), .CK(clock), .QN(n42) );
  DFF_X2 temp_yComputedVal_reg_6_ ( .D(n248), .CK(clock), .QN(n43) );
  DFF_X2 temp_yComputedVal_reg_5_ ( .D(n249), .CK(clock), .QN(n44) );
  DFF_X2 temp_yComputedVal_reg_4_ ( .D(n250), .CK(clock), .QN(n45) );
  DFF_X2 temp_yComputedVal_reg_3_ ( .D(n251), .CK(clock), .QN(n46) );
  DFF_X2 temp_yComputedVal_reg_2_ ( .D(n252), .CK(clock), .QN(n47) );
  DFF_X2 temp_yComputedVal_reg_1_ ( .D(n253), .CK(clock), .QN(n48) );
  DFF_X2 temp_yComputedVal_reg_0_ ( .D(n254), .CK(clock), .QN(n49) );
  DFF_X1 op_CPDoneFlag_reg ( .D(U11_Z_0), .CK(clock), .Q(op_CPDoneFlag) );
  OAI22_X2 U4 ( .A1(n154), .A2(n51), .B1(n53), .B2(n155), .ZN(n204) );
  NOR2_X2 U5 ( .A1(U16_DATA2_0), .A2(n156), .ZN(n155) );
  NAND3_X2 U7 ( .A1(n54), .A2(n52), .A3(U17_DATA2_0), .ZN(n157) );
  NAND2_X2 U8 ( .A1(n156), .A2(reset), .ZN(n154) );
  NAND2_X2 U9 ( .A1(n158), .A2(n55), .ZN(n206) );
  OAI22_X2 U11 ( .A1(n673), .A2(n2), .B1(n574), .B2(n106), .ZN(n207) );
  OAI22_X2 U12 ( .A1(n673), .A2(n3), .B1(n574), .B2(n107), .ZN(n208) );
  OAI22_X2 U13 ( .A1(n673), .A2(n4), .B1(n574), .B2(n108), .ZN(n209) );
  OAI22_X2 U14 ( .A1(n673), .A2(n5), .B1(n574), .B2(n109), .ZN(n210) );
  OAI22_X2 U22 ( .A1(n160), .A2(n13), .B1(n574), .B2(n117), .ZN(n218) );
  OAI22_X2 U23 ( .A1(n160), .A2(n14), .B1(n574), .B2(n118), .ZN(n219) );
  OAI22_X2 U24 ( .A1(n160), .A2(n15), .B1(n574), .B2(n119), .ZN(n220) );
  OAI22_X2 U25 ( .A1(n160), .A2(n16), .B1(n574), .B2(n120), .ZN(n221) );
  OAI22_X2 U26 ( .A1(n160), .A2(n17), .B1(n574), .B2(n121), .ZN(n222) );
  OAI22_X2 U27 ( .A1(n160), .A2(n18), .B1(n574), .B2(n122), .ZN(n223) );
  OAI22_X2 U28 ( .A1(n673), .A2(n19), .B1(n574), .B2(n123), .ZN(n224) );
  OAI22_X2 U29 ( .A1(n673), .A2(n20), .B1(n574), .B2(n124), .ZN(n225) );
  OAI22_X2 U30 ( .A1(n673), .A2(n21), .B1(n574), .B2(n125), .ZN(n226) );
  OAI22_X2 U31 ( .A1(n673), .A2(n22), .B1(n574), .B2(n126), .ZN(n227) );
  OAI22_X2 U32 ( .A1(n673), .A2(n23), .B1(n574), .B2(n127), .ZN(n228) );
  OAI22_X2 U33 ( .A1(n673), .A2(n24), .B1(n574), .B2(n128), .ZN(n229) );
  OAI22_X2 U34 ( .A1(n673), .A2(n25), .B1(n574), .B2(n129), .ZN(n230) );
  OAI22_X2 U35 ( .A1(n673), .A2(n26), .B1(n574), .B2(n130), .ZN(n231) );
  OAI22_X2 U36 ( .A1(n673), .A2(n27), .B1(n574), .B2(n131), .ZN(n232) );
  OAI22_X2 U37 ( .A1(n673), .A2(n28), .B1(n574), .B2(n132), .ZN(n233) );
  OAI22_X2 U38 ( .A1(n673), .A2(n29), .B1(n574), .B2(n133), .ZN(n234) );
  OAI22_X2 U39 ( .A1(n673), .A2(n30), .B1(n574), .B2(n134), .ZN(n235) );
  OAI22_X2 U40 ( .A1(n673), .A2(n31), .B1(n574), .B2(n135), .ZN(n236) );
  OAI22_X2 U41 ( .A1(n673), .A2(n32), .B1(n574), .B2(n136), .ZN(n237) );
  OAI22_X2 U42 ( .A1(n673), .A2(n33), .B1(n574), .B2(n137), .ZN(n238) );
  OAI22_X2 U43 ( .A1(n673), .A2(n34), .B1(n574), .B2(n138), .ZN(n239) );
  OAI22_X2 U44 ( .A1(n673), .A2(n35), .B1(n574), .B2(n139), .ZN(n240) );
  OAI22_X2 U45 ( .A1(n673), .A2(n36), .B1(n574), .B2(n140), .ZN(n241) );
  OAI22_X2 U46 ( .A1(n673), .A2(n37), .B1(n574), .B2(n141), .ZN(n242) );
  OAI22_X2 U47 ( .A1(n160), .A2(n38), .B1(n574), .B2(n142), .ZN(n243) );
  OAI22_X2 U48 ( .A1(n160), .A2(n39), .B1(n574), .B2(n143), .ZN(n244) );
  OAI22_X2 U49 ( .A1(n160), .A2(n40), .B1(n574), .B2(n144), .ZN(n245) );
  OAI22_X2 U50 ( .A1(n160), .A2(n41), .B1(n574), .B2(n145), .ZN(n246) );
  OAI22_X2 U51 ( .A1(n160), .A2(n42), .B1(n574), .B2(n146), .ZN(n247) );
  OAI22_X2 U52 ( .A1(n160), .A2(n43), .B1(n574), .B2(n147), .ZN(n248) );
  OAI22_X2 U53 ( .A1(n160), .A2(n44), .B1(n574), .B2(n148), .ZN(n249) );
  OAI22_X2 U54 ( .A1(n160), .A2(n45), .B1(n574), .B2(n149), .ZN(n250) );
  OAI22_X2 U55 ( .A1(n160), .A2(n46), .B1(n574), .B2(n150), .ZN(n251) );
  OAI22_X2 U56 ( .A1(n160), .A2(n47), .B1(n574), .B2(n151), .ZN(n252) );
  OAI22_X2 U57 ( .A1(n160), .A2(n48), .B1(n574), .B2(n152), .ZN(n253) );
  OAI22_X2 U58 ( .A1(n160), .A2(n49), .B1(n574), .B2(n153), .ZN(n254) );
  NAND2_X2 U59 ( .A1(n55), .A2(n50), .ZN(n160) );
  OAI22_X2 U60 ( .A1(n671), .A2(n96), .B1(n672), .B2(n40), .ZN(op_fpIn2[9]) );
  OAI22_X2 U61 ( .A1(n671), .A2(n97), .B1(n163), .B2(n41), .ZN(op_fpIn2[8]) );
  OAI22_X2 U62 ( .A1(n671), .A2(n98), .B1(n163), .B2(n42), .ZN(op_fpIn2[7]) );
  OAI22_X2 U63 ( .A1(n671), .A2(n99), .B1(n163), .B2(n43), .ZN(op_fpIn2[6]) );
  OAI22_X2 U64 ( .A1(n671), .A2(n100), .B1(n163), .B2(n44), .ZN(op_fpIn2[5])
         );
  OAI22_X2 U65 ( .A1(n671), .A2(n58), .B1(n163), .B2(n2), .ZN(op_fpIn2[47]) );
  OAI22_X2 U66 ( .A1(n671), .A2(n59), .B1(n163), .B2(n3), .ZN(op_fpIn2[46]) );
  OAI22_X2 U67 ( .A1(n671), .A2(n60), .B1(n163), .B2(n4), .ZN(op_fpIn2[45]) );
  OAI22_X2 U68 ( .A1(n671), .A2(n61), .B1(n163), .B2(n5), .ZN(op_fpIn2[44]) );
  OAI22_X2 U69 ( .A1(n671), .A2(n62), .B1(n163), .B2(n6), .ZN(op_fpIn2[43]) );
  OAI22_X2 U70 ( .A1(n671), .A2(n63), .B1(n163), .B2(n7), .ZN(op_fpIn2[42]) );
  OAI22_X2 U71 ( .A1(n671), .A2(n64), .B1(n163), .B2(n8), .ZN(op_fpIn2[41]) );
  OAI22_X2 U72 ( .A1(n671), .A2(n65), .B1(n163), .B2(n9), .ZN(op_fpIn2[40]) );
  OAI22_X2 U73 ( .A1(n671), .A2(n101), .B1(n163), .B2(n45), .ZN(op_fpIn2[4])
         );
  OAI22_X2 U74 ( .A1(n671), .A2(n66), .B1(n672), .B2(n10), .ZN(op_fpIn2[39])
         );
  OAI22_X2 U75 ( .A1(n671), .A2(n67), .B1(n672), .B2(n11), .ZN(op_fpIn2[38])
         );
  OAI22_X2 U76 ( .A1(n671), .A2(n68), .B1(n672), .B2(n12), .ZN(op_fpIn2[37])
         );
  OAI22_X2 U77 ( .A1(n671), .A2(n69), .B1(n672), .B2(n13), .ZN(op_fpIn2[36])
         );
  OAI22_X2 U78 ( .A1(n671), .A2(n70), .B1(n672), .B2(n14), .ZN(op_fpIn2[35])
         );
  OAI22_X2 U79 ( .A1(n671), .A2(n71), .B1(n672), .B2(n15), .ZN(op_fpIn2[34])
         );
  OAI22_X2 U80 ( .A1(n671), .A2(n72), .B1(n672), .B2(n16), .ZN(op_fpIn2[33])
         );
  OAI22_X2 U81 ( .A1(n671), .A2(n73), .B1(n672), .B2(n17), .ZN(op_fpIn2[32])
         );
  OAI22_X2 U82 ( .A1(n671), .A2(n74), .B1(n672), .B2(n18), .ZN(op_fpIn2[31])
         );
  OAI22_X2 U83 ( .A1(n671), .A2(n75), .B1(n672), .B2(n19), .ZN(op_fpIn2[30])
         );
  OAI22_X2 U84 ( .A1(n671), .A2(n102), .B1(n672), .B2(n46), .ZN(op_fpIn2[3])
         );
  OAI22_X2 U85 ( .A1(n671), .A2(n76), .B1(n672), .B2(n20), .ZN(op_fpIn2[29])
         );
  OAI22_X2 U86 ( .A1(n671), .A2(n77), .B1(n672), .B2(n21), .ZN(op_fpIn2[28])
         );
  OAI22_X2 U87 ( .A1(n671), .A2(n78), .B1(n672), .B2(n22), .ZN(op_fpIn2[27])
         );
  OAI22_X2 U88 ( .A1(n671), .A2(n79), .B1(n672), .B2(n23), .ZN(op_fpIn2[26])
         );
  OAI22_X2 U89 ( .A1(n671), .A2(n80), .B1(n672), .B2(n24), .ZN(op_fpIn2[25])
         );
  OAI22_X2 U90 ( .A1(n671), .A2(n81), .B1(n672), .B2(n25), .ZN(op_fpIn2[24])
         );
  OAI22_X2 U91 ( .A1(n671), .A2(n82), .B1(n672), .B2(n26), .ZN(op_fpIn2[23])
         );
  OAI22_X2 U92 ( .A1(n671), .A2(n83), .B1(n672), .B2(n27), .ZN(op_fpIn2[22])
         );
  OAI22_X2 U93 ( .A1(n671), .A2(n84), .B1(n672), .B2(n28), .ZN(op_fpIn2[21])
         );
  OAI22_X2 U94 ( .A1(n671), .A2(n85), .B1(n672), .B2(n29), .ZN(op_fpIn2[20])
         );
  OAI22_X2 U95 ( .A1(n671), .A2(n103), .B1(n672), .B2(n47), .ZN(op_fpIn2[2])
         );
  OAI22_X2 U96 ( .A1(n671), .A2(n86), .B1(n672), .B2(n30), .ZN(op_fpIn2[19])
         );
  OAI22_X2 U97 ( .A1(n671), .A2(n87), .B1(n672), .B2(n31), .ZN(op_fpIn2[18])
         );
  OAI22_X2 U98 ( .A1(n671), .A2(n88), .B1(n672), .B2(n32), .ZN(op_fpIn2[17])
         );
  OAI22_X2 U99 ( .A1(n671), .A2(n89), .B1(n672), .B2(n33), .ZN(op_fpIn2[16])
         );
  OAI22_X2 U100 ( .A1(n671), .A2(n90), .B1(n672), .B2(n34), .ZN(op_fpIn2[15])
         );
  OAI22_X2 U101 ( .A1(n671), .A2(n91), .B1(n672), .B2(n35), .ZN(op_fpIn2[14])
         );
  OAI22_X2 U102 ( .A1(n671), .A2(n92), .B1(n672), .B2(n36), .ZN(op_fpIn2[13])
         );
  OAI22_X2 U103 ( .A1(n671), .A2(n93), .B1(n672), .B2(n37), .ZN(op_fpIn2[12])
         );
  OAI22_X2 U104 ( .A1(n671), .A2(n94), .B1(n672), .B2(n38), .ZN(op_fpIn2[11])
         );
  OAI22_X2 U105 ( .A1(n671), .A2(n95), .B1(n672), .B2(n39), .ZN(op_fpIn2[10])
         );
  OAI22_X2 U106 ( .A1(n671), .A2(n104), .B1(n672), .B2(n48), .ZN(op_fpIn2[1])
         );
  OAI22_X2 U107 ( .A1(n671), .A2(n105), .B1(n163), .B2(n49), .ZN(op_fpIn2[0])
         );
  NOR2_X2 U108 ( .A1(n57), .A2(n164), .ZN(n163) );
  NOR2_X2 U109 ( .A1(n52), .A2(n156), .ZN(U11_Z_0) );
  NAND2_X2 U110 ( .A1(n159), .A2(n55), .ZN(n156) );
  NAND2_X2 U111 ( .A1(executeEnableBit), .A2(reset), .ZN(n162) );
  NOR2_X2 U112 ( .A1(n165), .A2(n164), .ZN(n159) );
  NOR4_X2 U113 ( .A1(n166), .A2(n167), .A3(n168), .A4(n169), .ZN(n164) );
  NAND4_X2 U114 ( .A1(n170), .A2(n171), .A3(n172), .A4(n173), .ZN(n169) );
  NOR3_X2 U115 ( .A1(yInVal1[3]), .A2(yInVal1[41]), .A3(yInVal1[40]), .ZN(n173) );
  NOR3_X2 U116 ( .A1(yInVal1[37]), .A2(yInVal1[39]), .A3(yInVal1[38]), .ZN(
        n172) );
  NOR3_X2 U117 ( .A1(yInVal1[34]), .A2(yInVal1[36]), .A3(yInVal1[35]), .ZN(
        n171) );
  NOR3_X2 U118 ( .A1(yInVal1[31]), .A2(yInVal1[33]), .A3(yInVal1[32]), .ZN(
        n170) );
  NAND4_X2 U119 ( .A1(n174), .A2(n175), .A3(n176), .A4(n177), .ZN(n168) );
  NOR3_X2 U120 ( .A1(yInVal1[7]), .A2(yInVal1[9]), .A3(yInVal1[8]), .ZN(n177)
         );
  NOR3_X2 U121 ( .A1(yInVal1[4]), .A2(yInVal1[6]), .A3(yInVal1[5]), .ZN(n176)
         );
  NOR3_X2 U122 ( .A1(yInVal1[45]), .A2(yInVal1[47]), .A3(yInVal1[46]), .ZN(
        n175) );
  NOR3_X2 U123 ( .A1(yInVal1[42]), .A2(yInVal1[44]), .A3(yInVal1[43]), .ZN(
        n174) );
  NAND4_X2 U124 ( .A1(n178), .A2(n179), .A3(n180), .A4(n181), .ZN(n167) );
  NOR3_X2 U125 ( .A1(yInVal1[18]), .A2(yInVal1[1]), .A3(yInVal1[19]), .ZN(n181) );
  NOR3_X2 U126 ( .A1(yInVal1[15]), .A2(yInVal1[17]), .A3(yInVal1[16]), .ZN(
        n180) );
  NOR3_X2 U127 ( .A1(yInVal1[12]), .A2(yInVal1[14]), .A3(yInVal1[13]), .ZN(
        n179) );
  NOR3_X2 U128 ( .A1(yInVal1[0]), .A2(yInVal1[11]), .A3(yInVal1[10]), .ZN(n178) );
  NAND4_X2 U129 ( .A1(n182), .A2(n183), .A3(n184), .A4(n185), .ZN(n166) );
  NOR3_X2 U130 ( .A1(yInVal1[29]), .A2(yInVal1[30]), .A3(yInVal1[2]), .ZN(n185) );
  NOR3_X2 U131 ( .A1(yInVal1[26]), .A2(yInVal1[28]), .A3(yInVal1[27]), .ZN(
        n184) );
  NOR3_X2 U132 ( .A1(yInVal1[23]), .A2(yInVal1[25]), .A3(yInVal1[24]), .ZN(
        n183) );
  NOR3_X2 U133 ( .A1(yInVal1[20]), .A2(yInVal1[22]), .A3(yInVal1[21]), .ZN(
        n182) );
  NAND2_X2 U134 ( .A1(n186), .A2(n187), .ZN(n165) );
  NOR4_X2 U135 ( .A1(n188), .A2(n189), .A3(n190), .A4(n191), .ZN(n187) );
  NAND4_X2 U136 ( .A1(n74), .A2(n73), .A3(n75), .A4(n192), .ZN(n191) );
  NOR3_X2 U137 ( .A1(yInVal2[33]), .A2(yInVal2[35]), .A3(yInVal2[34]), .ZN(
        n192) );
  NAND4_X2 U138 ( .A1(n68), .A2(n67), .A3(n69), .A4(n193), .ZN(n190) );
  NOR3_X2 U139 ( .A1(yInVal2[39]), .A2(yInVal2[40]), .A3(yInVal2[4]), .ZN(n193) );
  NAND4_X2 U140 ( .A1(n63), .A2(n62), .A3(n64), .A4(n194), .ZN(n189) );
  NOR3_X2 U141 ( .A1(yInVal2[44]), .A2(yInVal2[46]), .A3(yInVal2[45]), .ZN(
        n194) );
  NAND4_X2 U142 ( .A1(n100), .A2(n99), .A3(n58), .A4(n195), .ZN(n188) );
  NOR3_X2 U143 ( .A1(yInVal2[7]), .A2(yInVal2[9]), .A3(yInVal2[8]), .ZN(n195)
         );
  NOR4_X2 U144 ( .A1(n196), .A2(n197), .A3(n198), .A4(n199), .ZN(n186) );
  NAND4_X2 U145 ( .A1(n104), .A2(n95), .A3(n105), .A4(n200), .ZN(n199) );
  NOR3_X2 U146 ( .A1(yInVal2[11]), .A2(yInVal2[13]), .A3(yInVal2[12]), .ZN(
        n200) );
  NAND4_X2 U147 ( .A1(n90), .A2(n89), .A3(n91), .A4(n201), .ZN(n198) );
  NOR3_X2 U148 ( .A1(yInVal2[17]), .A2(yInVal2[19]), .A3(yInVal2[18]), .ZN(
        n201) );
  NAND4_X2 U149 ( .A1(n85), .A2(n84), .A3(n103), .A4(n202), .ZN(n197) );
  NOR3_X2 U150 ( .A1(yInVal2[22]), .A2(yInVal2[24]), .A3(yInVal2[23]), .ZN(
        n202) );
  NAND4_X2 U151 ( .A1(n79), .A2(n78), .A3(n80), .A4(n203), .ZN(n196) );
  NOR3_X2 U152 ( .A1(yInVal2[28]), .A2(yInVal2[3]), .A3(yInVal2[29]), .ZN(n203) );
  INV_X4 U153 ( .A(n154), .ZN(n53) );
  INV_X4 U154 ( .A(n156), .ZN(n54) );
  INV_X4 U155 ( .A(n162), .ZN(n55) );
  INV_X4 U157 ( .A(n165), .ZN(n57) );
  INV_X4 U158 ( .A(yInVal2[47]), .ZN(n58) );
  INV_X4 U159 ( .A(yInVal2[46]), .ZN(n59) );
  INV_X4 U160 ( .A(yInVal2[45]), .ZN(n60) );
  INV_X4 U161 ( .A(yInVal2[44]), .ZN(n61) );
  INV_X4 U162 ( .A(yInVal2[43]), .ZN(n62) );
  INV_X4 U163 ( .A(yInVal2[42]), .ZN(n63) );
  INV_X4 U164 ( .A(yInVal2[41]), .ZN(n64) );
  INV_X4 U165 ( .A(yInVal2[40]), .ZN(n65) );
  INV_X4 U166 ( .A(yInVal2[39]), .ZN(n66) );
  INV_X4 U167 ( .A(yInVal2[38]), .ZN(n67) );
  INV_X4 U168 ( .A(yInVal2[37]), .ZN(n68) );
  INV_X4 U169 ( .A(yInVal2[36]), .ZN(n69) );
  INV_X4 U170 ( .A(yInVal2[35]), .ZN(n70) );
  INV_X4 U171 ( .A(yInVal2[34]), .ZN(n71) );
  INV_X4 U172 ( .A(yInVal2[33]), .ZN(n72) );
  INV_X4 U173 ( .A(yInVal2[32]), .ZN(n73) );
  INV_X4 U174 ( .A(yInVal2[31]), .ZN(n74) );
  INV_X4 U175 ( .A(yInVal2[30]), .ZN(n75) );
  INV_X4 U176 ( .A(yInVal2[29]), .ZN(n76) );
  INV_X4 U177 ( .A(yInVal2[28]), .ZN(n77) );
  INV_X4 U178 ( .A(yInVal2[27]), .ZN(n78) );
  INV_X4 U179 ( .A(yInVal2[26]), .ZN(n79) );
  INV_X4 U180 ( .A(yInVal2[25]), .ZN(n80) );
  INV_X4 U181 ( .A(yInVal2[24]), .ZN(n81) );
  INV_X4 U182 ( .A(yInVal2[23]), .ZN(n82) );
  INV_X4 U183 ( .A(yInVal2[22]), .ZN(n83) );
  INV_X4 U184 ( .A(yInVal2[21]), .ZN(n84) );
  INV_X4 U185 ( .A(yInVal2[20]), .ZN(n85) );
  INV_X4 U186 ( .A(yInVal2[19]), .ZN(n86) );
  INV_X4 U187 ( .A(yInVal2[18]), .ZN(n87) );
  INV_X4 U188 ( .A(yInVal2[17]), .ZN(n88) );
  INV_X4 U189 ( .A(yInVal2[16]), .ZN(n89) );
  INV_X4 U190 ( .A(yInVal2[15]), .ZN(n90) );
  INV_X4 U191 ( .A(yInVal2[14]), .ZN(n91) );
  INV_X4 U192 ( .A(yInVal2[13]), .ZN(n92) );
  INV_X4 U193 ( .A(yInVal2[12]), .ZN(n93) );
  INV_X4 U194 ( .A(yInVal2[11]), .ZN(n94) );
  INV_X4 U195 ( .A(yInVal2[10]), .ZN(n95) );
  INV_X4 U196 ( .A(yInVal2[9]), .ZN(n96) );
  INV_X4 U197 ( .A(yInVal2[8]), .ZN(n97) );
  INV_X4 U198 ( .A(yInVal2[7]), .ZN(n98) );
  INV_X4 U199 ( .A(yInVal2[6]), .ZN(n99) );
  INV_X4 U200 ( .A(yInVal2[5]), .ZN(n100) );
  INV_X4 U201 ( .A(yInVal2[4]), .ZN(n101) );
  INV_X4 U202 ( .A(yInVal2[3]), .ZN(n102) );
  INV_X4 U203 ( .A(yInVal2[2]), .ZN(n103) );
  INV_X4 U204 ( .A(yInVal2[1]), .ZN(n104) );
  INV_X4 U205 ( .A(yInVal2[0]), .ZN(n105) );
  INV_X4 U206 ( .A(in_fpOut[47]), .ZN(n106) );
  INV_X4 U207 ( .A(in_fpOut[46]), .ZN(n107) );
  INV_X4 U208 ( .A(in_fpOut[45]), .ZN(n108) );
  INV_X4 U209 ( .A(in_fpOut[44]), .ZN(n109) );
  INV_X4 U210 ( .A(in_fpOut[43]), .ZN(n110) );
  INV_X4 U211 ( .A(in_fpOut[42]), .ZN(n111) );
  INV_X4 U212 ( .A(in_fpOut[41]), .ZN(n112) );
  INV_X4 U213 ( .A(in_fpOut[40]), .ZN(n113) );
  INV_X4 U214 ( .A(in_fpOut[39]), .ZN(n114) );
  INV_X4 U215 ( .A(in_fpOut[38]), .ZN(n115) );
  INV_X4 U216 ( .A(in_fpOut[37]), .ZN(n116) );
  INV_X4 U217 ( .A(in_fpOut[36]), .ZN(n117) );
  INV_X4 U218 ( .A(in_fpOut[35]), .ZN(n118) );
  INV_X4 U219 ( .A(in_fpOut[34]), .ZN(n119) );
  INV_X4 U220 ( .A(in_fpOut[33]), .ZN(n120) );
  INV_X4 U221 ( .A(in_fpOut[32]), .ZN(n121) );
  INV_X4 U222 ( .A(in_fpOut[31]), .ZN(n122) );
  INV_X4 U223 ( .A(in_fpOut[30]), .ZN(n123) );
  INV_X4 U224 ( .A(in_fpOut[29]), .ZN(n124) );
  INV_X4 U225 ( .A(in_fpOut[28]), .ZN(n125) );
  INV_X4 U226 ( .A(in_fpOut[27]), .ZN(n126) );
  INV_X4 U227 ( .A(in_fpOut[26]), .ZN(n127) );
  INV_X4 U228 ( .A(in_fpOut[25]), .ZN(n128) );
  INV_X4 U229 ( .A(in_fpOut[24]), .ZN(n129) );
  INV_X4 U230 ( .A(in_fpOut[23]), .ZN(n130) );
  INV_X4 U231 ( .A(in_fpOut[22]), .ZN(n131) );
  INV_X4 U232 ( .A(in_fpOut[21]), .ZN(n132) );
  INV_X4 U233 ( .A(in_fpOut[20]), .ZN(n133) );
  INV_X4 U234 ( .A(in_fpOut[19]), .ZN(n134) );
  INV_X4 U235 ( .A(in_fpOut[18]), .ZN(n135) );
  INV_X4 U236 ( .A(in_fpOut[17]), .ZN(n136) );
  INV_X4 U237 ( .A(in_fpOut[16]), .ZN(n137) );
  INV_X4 U238 ( .A(in_fpOut[15]), .ZN(n138) );
  INV_X4 U239 ( .A(in_fpOut[14]), .ZN(n139) );
  INV_X4 U240 ( .A(in_fpOut[13]), .ZN(n140) );
  INV_X4 U241 ( .A(in_fpOut[12]), .ZN(n141) );
  INV_X4 U242 ( .A(in_fpOut[11]), .ZN(n142) );
  INV_X4 U243 ( .A(in_fpOut[10]), .ZN(n143) );
  INV_X4 U244 ( .A(in_fpOut[9]), .ZN(n144) );
  INV_X4 U245 ( .A(in_fpOut[8]), .ZN(n145) );
  INV_X4 U246 ( .A(in_fpOut[7]), .ZN(n146) );
  INV_X4 U247 ( .A(in_fpOut[6]), .ZN(n147) );
  INV_X4 U248 ( .A(in_fpOut[5]), .ZN(n148) );
  INV_X4 U249 ( .A(in_fpOut[4]), .ZN(n149) );
  INV_X4 U250 ( .A(in_fpOut[3]), .ZN(n150) );
  INV_X4 U251 ( .A(in_fpOut[2]), .ZN(n151) );
  INV_X4 U252 ( .A(in_fpOut[1]), .ZN(n152) );
  INV_X4 U253 ( .A(in_fpOut[0]), .ZN(n153) );
  DFF_X2 temp_nextMode_reg ( .D(n206), .CK(clock), .Q(op_fpMode) );
  DFF_X2 temp_count_for_CPDoneFlag_reg_0_ ( .D(n205), .CK(clock), .Q(
        U16_DATA2_0), .QN(n52) );
  DFF_X2 temp_count_for_CPDoneFlag_reg_1_ ( .D(n204), .CK(clock), .Q(
        U17_DATA2_0), .QN(n51) );
  OR3_X4 U6 ( .A1(op_DoneFlag), .A2(n162), .A3(n50), .ZN(n574) );
  INV_X4 U156 ( .A(n671), .ZN(n672) );
  INV_X4 U254 ( .A(n674), .ZN(n673) );
  BUF_X4 U255 ( .A(in_fpOut[0]), .Z(op_yWriteVal[0]) );
  BUF_X4 U256 ( .A(in_fpOut[1]), .Z(op_yWriteVal[1]) );
  BUF_X4 U257 ( .A(in_fpOut[2]), .Z(op_yWriteVal[2]) );
  BUF_X4 U258 ( .A(in_fpOut[3]), .Z(op_yWriteVal[3]) );
  BUF_X4 U259 ( .A(in_fpOut[4]), .Z(op_yWriteVal[4]) );
  BUF_X4 U260 ( .A(in_fpOut[5]), .Z(op_yWriteVal[5]) );
  BUF_X4 U261 ( .A(in_fpOut[6]), .Z(op_yWriteVal[6]) );
  BUF_X4 U262 ( .A(in_fpOut[7]), .Z(op_yWriteVal[7]) );
  BUF_X4 U263 ( .A(in_fpOut[8]), .Z(op_yWriteVal[8]) );
  BUF_X4 U264 ( .A(in_fpOut[9]), .Z(op_yWriteVal[9]) );
  BUF_X4 U265 ( .A(in_fpOut[10]), .Z(op_yWriteVal[10]) );
  BUF_X4 U266 ( .A(in_fpOut[11]), .Z(op_yWriteVal[11]) );
  BUF_X4 U267 ( .A(in_fpOut[12]), .Z(op_yWriteVal[12]) );
  BUF_X4 U268 ( .A(in_fpOut[13]), .Z(op_yWriteVal[13]) );
  BUF_X4 U269 ( .A(in_fpOut[14]), .Z(op_yWriteVal[14]) );
  BUF_X4 U270 ( .A(in_fpOut[15]), .Z(op_yWriteVal[15]) );
  BUF_X4 U271 ( .A(in_fpOut[16]), .Z(op_yWriteVal[16]) );
  BUF_X4 U272 ( .A(in_fpOut[17]), .Z(op_yWriteVal[17]) );
  BUF_X4 U273 ( .A(in_fpOut[18]), .Z(op_yWriteVal[18]) );
  BUF_X4 U274 ( .A(in_fpOut[19]), .Z(op_yWriteVal[19]) );
  BUF_X4 U275 ( .A(in_fpOut[20]), .Z(op_yWriteVal[20]) );
  BUF_X4 U276 ( .A(in_fpOut[21]), .Z(op_yWriteVal[21]) );
  BUF_X4 U277 ( .A(in_fpOut[22]), .Z(op_yWriteVal[22]) );
  BUF_X4 U278 ( .A(in_fpOut[23]), .Z(op_yWriteVal[23]) );
  BUF_X4 U279 ( .A(in_fpOut[24]), .Z(op_yWriteVal[24]) );
  INV_X4 U280 ( .A(n160), .ZN(n674) );
  OAI21_X2 U281 ( .B1(n52), .B2(n154), .A(n157), .ZN(n205) );
  AOI21_X1 U282 ( .B1(op_fpMode), .B2(n671), .A(n159), .ZN(n158) );
  BUF_X4 U283 ( .A(yInVal1[0]), .Z(op_fpIn1[0]) );
  BUF_X4 U284 ( .A(yInVal1[1]), .Z(op_fpIn1[1]) );
  BUF_X4 U285 ( .A(yInVal1[2]), .Z(op_fpIn1[2]) );
  BUF_X4 U286 ( .A(yInVal1[3]), .Z(op_fpIn1[3]) );
  BUF_X4 U287 ( .A(yInVal1[4]), .Z(op_fpIn1[4]) );
  BUF_X4 U288 ( .A(yInVal1[5]), .Z(op_fpIn1[5]) );
  BUF_X4 U289 ( .A(yInVal1[6]), .Z(op_fpIn1[6]) );
  BUF_X4 U290 ( .A(yInVal1[7]), .Z(op_fpIn1[7]) );
  BUF_X4 U291 ( .A(yInVal1[8]), .Z(op_fpIn1[8]) );
  BUF_X4 U292 ( .A(yInVal1[9]), .Z(op_fpIn1[9]) );
  BUF_X4 U293 ( .A(yInVal1[10]), .Z(op_fpIn1[10]) );
  BUF_X4 U294 ( .A(yInVal1[11]), .Z(op_fpIn1[11]) );
  BUF_X4 U295 ( .A(yInVal1[12]), .Z(op_fpIn1[12]) );
  BUF_X4 U296 ( .A(yInVal1[13]), .Z(op_fpIn1[13]) );
  BUF_X4 U297 ( .A(yInVal1[14]), .Z(op_fpIn1[14]) );
  BUF_X4 U298 ( .A(yInVal1[15]), .Z(op_fpIn1[15]) );
  BUF_X4 U299 ( .A(yInVal1[16]), .Z(op_fpIn1[16]) );
  BUF_X4 U300 ( .A(yInVal1[17]), .Z(op_fpIn1[17]) );
  BUF_X4 U301 ( .A(yInVal1[18]), .Z(op_fpIn1[18]) );
  BUF_X4 U302 ( .A(yInVal1[19]), .Z(op_fpIn1[19]) );
  BUF_X4 U303 ( .A(yInVal1[20]), .Z(op_fpIn1[20]) );
  BUF_X4 U304 ( .A(yInVal1[21]), .Z(op_fpIn1[21]) );
  BUF_X4 U305 ( .A(yInVal1[22]), .Z(op_fpIn1[22]) );
  BUF_X4 U306 ( .A(yInVal1[23]), .Z(op_fpIn1[23]) );
  BUF_X4 U307 ( .A(yInVal1[24]), .Z(op_fpIn1[24]) );
  BUF_X4 U308 ( .A(yInVal1[25]), .Z(op_fpIn1[25]) );
  BUF_X4 U309 ( .A(yInVal1[26]), .Z(op_fpIn1[26]) );
  BUF_X4 U310 ( .A(yInVal1[27]), .Z(op_fpIn1[27]) );
  BUF_X4 U311 ( .A(yInVal1[28]), .Z(op_fpIn1[28]) );
  BUF_X4 U312 ( .A(yInVal1[29]), .Z(op_fpIn1[29]) );
  BUF_X4 U313 ( .A(yInVal1[30]), .Z(op_fpIn1[30]) );
  BUF_X4 U314 ( .A(yInVal1[31]), .Z(op_fpIn1[31]) );
  BUF_X4 U315 ( .A(yInVal1[32]), .Z(op_fpIn1[32]) );
  BUF_X4 U316 ( .A(yInVal1[33]), .Z(op_fpIn1[33]) );
  BUF_X4 U317 ( .A(yInVal1[34]), .Z(op_fpIn1[34]) );
  BUF_X4 U318 ( .A(yInVal1[35]), .Z(op_fpIn1[35]) );
  BUF_X4 U319 ( .A(yInVal1[36]), .Z(op_fpIn1[36]) );
  BUF_X4 U320 ( .A(yInVal1[37]), .Z(op_fpIn1[37]) );
  BUF_X4 U321 ( .A(yInVal1[38]), .Z(op_fpIn1[38]) );
  BUF_X4 U322 ( .A(yInVal1[39]), .Z(op_fpIn1[39]) );
  BUF_X4 U323 ( .A(yInVal1[40]), .Z(op_fpIn1[40]) );
  BUF_X4 U324 ( .A(yInVal1[41]), .Z(op_fpIn1[41]) );
  BUF_X4 U325 ( .A(yInVal1[42]), .Z(op_fpIn1[42]) );
  BUF_X4 U326 ( .A(yInVal1[43]), .Z(op_fpIn1[43]) );
  BUF_X4 U327 ( .A(yInVal1[44]), .Z(op_fpIn1[44]) );
  BUF_X4 U328 ( .A(yInVal1[45]), .Z(op_fpIn1[45]) );
  BUF_X4 U329 ( .A(yInVal1[46]), .Z(op_fpIn1[46]) );
  BUF_X4 U330 ( .A(yInVal1[47]), .Z(op_fpIn1[47]) );
  BUF_X4 U331 ( .A(in_fpOut[47]), .Z(op_yWriteVal[47]) );
  BUF_X4 U332 ( .A(in_fpOut[46]), .Z(op_yWriteVal[46]) );
  BUF_X4 U333 ( .A(in_fpOut[45]), .Z(op_yWriteVal[45]) );
  BUF_X4 U334 ( .A(in_fpOut[44]), .Z(op_yWriteVal[44]) );
  BUF_X4 U335 ( .A(in_fpOut[43]), .Z(op_yWriteVal[43]) );
  BUF_X4 U336 ( .A(in_fpOut[42]), .Z(op_yWriteVal[42]) );
  BUF_X4 U337 ( .A(in_fpOut[41]), .Z(op_yWriteVal[41]) );
  BUF_X4 U338 ( .A(in_fpOut[40]), .Z(op_yWriteVal[40]) );
  BUF_X4 U339 ( .A(in_fpOut[39]), .Z(op_yWriteVal[39]) );
  BUF_X4 U340 ( .A(in_fpOut[38]), .Z(op_yWriteVal[38]) );
  BUF_X4 U341 ( .A(in_fpOut[37]), .Z(op_yWriteVal[37]) );
  BUF_X4 U342 ( .A(in_fpOut[36]), .Z(op_yWriteVal[36]) );
  BUF_X4 U343 ( .A(in_fpOut[35]), .Z(op_yWriteVal[35]) );
  BUF_X4 U344 ( .A(in_fpOut[34]), .Z(op_yWriteVal[34]) );
  BUF_X4 U345 ( .A(in_fpOut[33]), .Z(op_yWriteVal[33]) );
  BUF_X4 U346 ( .A(in_fpOut[32]), .Z(op_yWriteVal[32]) );
  BUF_X4 U347 ( .A(in_fpOut[31]), .Z(op_yWriteVal[31]) );
  BUF_X4 U348 ( .A(in_fpOut[30]), .Z(op_yWriteVal[30]) );
  BUF_X4 U349 ( .A(in_fpOut[29]), .Z(op_yWriteVal[29]) );
  BUF_X4 U350 ( .A(in_fpOut[28]), .Z(op_yWriteVal[28]) );
  BUF_X4 U351 ( .A(in_fpOut[27]), .Z(op_yWriteVal[27]) );
  BUF_X4 U352 ( .A(in_fpOut[26]), .Z(op_yWriteVal[26]) );
  BUF_X4 U353 ( .A(in_fpOut[25]), .Z(op_yWriteVal[25]) );
  OAI22_X1 U10 ( .A1(n160), .A2(n6), .B1(n574), .B2(n110), .ZN(n211) );
  OAI22_X1 U15 ( .A1(n160), .A2(n7), .B1(n574), .B2(n111), .ZN(n212) );
  OAI22_X1 U16 ( .A1(n160), .A2(n8), .B1(n574), .B2(n112), .ZN(n213) );
  OAI22_X1 U17 ( .A1(n160), .A2(n9), .B1(n574), .B2(n113), .ZN(n214) );
  OAI22_X1 U18 ( .A1(n160), .A2(n10), .B1(n574), .B2(n114), .ZN(n215) );
  OAI22_X1 U19 ( .A1(n160), .A2(n11), .B1(n574), .B2(n115), .ZN(n216) );
  OAI22_X1 U20 ( .A1(n160), .A2(n12), .B1(n574), .B2(n116), .ZN(n217) );
  INV_X8 U21 ( .A(n163), .ZN(n671) );
endmodule


module updateY_control ( clock, reset, exModDone, chng_row, chng_col, 
        chng_real, chng_img, dpModDoneFlag, ymem_data1, ymem_data2, filt_EN, 
        yMemDataReadyNextCycle, yAddrIn1, yAddrIn2, op_y_row, op_yVal1, 
        op_yVal2, op_EX_EN, op_DataEN, op_yAddrDiag, op_yAddrNonDiag, 
        op_oneHotDiag, op_oneHotNonDiag );
  input [15:0] chng_row;
  input [15:0] chng_col;
  input [23:0] chng_real;
  input [23:0] chng_img;
  input [255:0] ymem_data1;
  input [255:0] ymem_data2;
  input [10:0] yAddrIn1;
  input [10:0] yAddrIn2;
  output [15:0] op_y_row;
  output [47:0] op_yVal1;
  output [47:0] op_yVal2;
  output [10:0] op_yAddrDiag;
  output [10:0] op_yAddrNonDiag;
  output [3:0] op_oneHotDiag;
  output [3:0] op_oneHotNonDiag;
  input clock, reset, exModDone, dpModDoneFlag, filt_EN,
         yMemDataReadyNextCycle;
  output op_EX_EN, op_DataEN;
  wire   U95_Z_0, U95_Z_1, U95_Z_2, U94_Z_0, U94_Z_1, U94_Z_2, U94_Z_3,
         U94_Z_4, U94_Z_5, U94_Z_6, U94_Z_7, U94_Z_8, U94_Z_9, U94_Z_10,
         U94_Z_11, U94_Z_12, U94_Z_13, U94_Z_14, U94_Z_15, U94_Z_16, U94_Z_17,
         U94_Z_18, U94_Z_19, U94_Z_20, U94_Z_21, U94_Z_22, U94_Z_23, U94_Z_24,
         U94_Z_25, U94_Z_26, U94_Z_27, U94_Z_28, U94_Z_29, U94_Z_30, U94_Z_31,
         U94_Z_32, U94_Z_33, U94_Z_34, U94_Z_35, U94_Z_36, U94_Z_37, U94_Z_38,
         U94_Z_39, U94_Z_40, U94_Z_41, U94_Z_42, U94_Z_43, U94_Z_44, U94_Z_45,
         U94_Z_46, U94_Z_47, U93_Z_0, U93_Z_1, U93_Z_2, U93_Z_3, U93_Z_4,
         U93_Z_5, U93_Z_6, U93_Z_7, U93_Z_8, U93_Z_9, U93_Z_10, U93_Z_11,
         U93_Z_12, U93_Z_13, U93_Z_14, U93_Z_15, U93_Z_16, U93_Z_17, U93_Z_18,
         U93_Z_19, U93_Z_20, U93_Z_21, U93_Z_22, U93_Z_23, U93_Z_24, U93_Z_25,
         U93_Z_26, U93_Z_27, U93_Z_28, U93_Z_29, U93_Z_30, U93_Z_31, U93_Z_32,
         U93_Z_33, U93_Z_34, U93_Z_35, U93_Z_36, U93_Z_37, U93_Z_38, U93_Z_39,
         U93_Z_40, U93_Z_41, U93_Z_42, U93_Z_43, U93_Z_44, U93_Z_45, U93_Z_46,
         U93_Z_47, U92_Z_0, U91_Z_0, U91_Z_1, U91_Z_2, U91_Z_3, U91_Z_4,
         U91_Z_5, U91_Z_6, U91_Z_7, U91_Z_8, U91_Z_9, U91_Z_10, U91_Z_11,
         U91_Z_12, U91_Z_13, U91_Z_14, U91_Z_15, U90_Z_0, U72_DATA1_0,
         U72_DATA1_1, U72_DATA1_2, U72_DATA1_3, U72_DATA1_4, U72_DATA1_5,
         U72_DATA1_6, U72_DATA1_7, U72_DATA1_8, U72_DATA1_9, U72_DATA1_10,
         U72_DATA1_11, U72_DATA1_12, U72_DATA1_13, U72_DATA1_14, U72_DATA1_15,
         U72_DATA1_16, U72_DATA1_17, U72_DATA1_18, U72_DATA1_19, U72_DATA1_20,
         U72_DATA1_21, U72_DATA1_22, U72_DATA1_23, U72_DATA1_24, U72_DATA1_25,
         U72_DATA1_26, U72_DATA1_27, U72_DATA1_28, U72_DATA1_29, U72_DATA1_30,
         U72_DATA1_31, U72_DATA1_32, U72_DATA1_33, U72_DATA1_34, U72_DATA1_35,
         U72_DATA1_36, U72_DATA1_37, U72_DATA1_38, U72_DATA1_39, U72_DATA1_40,
         U72_DATA1_41, U72_DATA1_42, U72_DATA1_43, U72_DATA1_44, U72_DATA1_45,
         U72_DATA1_46, U72_DATA1_47, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n105, n107, n109, n110, n111, n112,
         n113, n115, n116, n117, n118, n120, n121, n122, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n141, n145, n146, n149, n150, n151, n152, n153, n154,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n782, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n801, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n831, n832, n834, n835,
         n837, n838, n839, n840, n841, n843, n844, n845, n846, n849, n850,
         n851, n852, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1807,
         n1808, n1810, n1811, n1813, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309;
  wire   [2372:2370] n;

  DFF_X1 op_oneHotNonDiag_reg_1_ ( .D(n2628), .CK(clock), .Q(
        op_oneHotNonDiag[1]) );
  DFF_X1 op_oneHotNonDiag_reg_0_ ( .D(n1), .CK(clock), .Q(op_oneHotNonDiag[0])
         );
  DFF_X1 op_oneHotNonDiag_reg_2_ ( .D(n2629), .CK(clock), .Q(
        op_oneHotNonDiag[2]) );
  DFF_X1 op_oneHotNonDiag_reg_3_ ( .D(n2630), .CK(clock), .Q(
        op_oneHotNonDiag[3]) );
  DFF_X1 temp_yVal_reg_0_ ( .D(n2631), .CK(clock), .Q(U72_DATA1_0), .QN(n58)
         );
  DFF_X1 temp_yVal_reg_1_ ( .D(n2632), .CK(clock), .Q(U72_DATA1_1), .QN(n57)
         );
  DFF_X1 temp_yVal_reg_2_ ( .D(n2633), .CK(clock), .Q(U72_DATA1_2), .QN(n56)
         );
  DFF_X1 temp_yVal_reg_3_ ( .D(n2634), .CK(clock), .Q(U72_DATA1_3), .QN(n55)
         );
  DFF_X1 temp_yVal_reg_4_ ( .D(n2635), .CK(clock), .Q(U72_DATA1_4), .QN(n54)
         );
  DFF_X1 temp_yVal_reg_5_ ( .D(n2636), .CK(clock), .Q(U72_DATA1_5), .QN(n53)
         );
  DFF_X1 temp_yVal_reg_6_ ( .D(n2637), .CK(clock), .Q(U72_DATA1_6), .QN(n52)
         );
  DFF_X1 temp_yVal_reg_7_ ( .D(n2638), .CK(clock), .Q(U72_DATA1_7), .QN(n51)
         );
  DFF_X1 temp_yVal_reg_8_ ( .D(n2639), .CK(clock), .Q(U72_DATA1_8), .QN(n50)
         );
  DFF_X1 temp_yVal_reg_9_ ( .D(n2640), .CK(clock), .Q(U72_DATA1_9), .QN(n49)
         );
  DFF_X1 temp_yVal_reg_10_ ( .D(n2641), .CK(clock), .Q(U72_DATA1_10), .QN(n48)
         );
  DFF_X1 temp_yVal_reg_11_ ( .D(n2642), .CK(clock), .Q(U72_DATA1_11), .QN(n47)
         );
  DFF_X1 temp_yVal_reg_12_ ( .D(n2643), .CK(clock), .Q(U72_DATA1_12), .QN(n46)
         );
  DFF_X1 temp_yVal_reg_13_ ( .D(n2644), .CK(clock), .Q(U72_DATA1_13), .QN(n45)
         );
  DFF_X1 temp_yVal_reg_14_ ( .D(n2645), .CK(clock), .Q(U72_DATA1_14), .QN(n44)
         );
  DFF_X1 temp_yVal_reg_15_ ( .D(n2646), .CK(clock), .Q(U72_DATA1_15), .QN(n43)
         );
  DFF_X1 temp_yVal_reg_16_ ( .D(n2647), .CK(clock), .Q(U72_DATA1_16), .QN(n42)
         );
  DFF_X1 temp_yVal_reg_17_ ( .D(n2648), .CK(clock), .Q(U72_DATA1_17), .QN(n41)
         );
  DFF_X1 temp_yVal_reg_18_ ( .D(n2649), .CK(clock), .Q(U72_DATA1_18), .QN(n40)
         );
  DFF_X1 temp_yVal_reg_19_ ( .D(n2650), .CK(clock), .Q(U72_DATA1_19), .QN(n39)
         );
  DFF_X1 temp_yVal_reg_20_ ( .D(n2651), .CK(clock), .Q(U72_DATA1_20), .QN(n38)
         );
  DFF_X1 temp_yVal_reg_21_ ( .D(n2652), .CK(clock), .Q(U72_DATA1_21), .QN(n37)
         );
  DFF_X1 temp_yVal_reg_22_ ( .D(n2653), .CK(clock), .Q(U72_DATA1_22), .QN(n36)
         );
  DFF_X1 temp_yVal_reg_23_ ( .D(n2654), .CK(clock), .Q(U72_DATA1_23), .QN(n35)
         );
  DFF_X1 temp_yVal_reg_24_ ( .D(n2655), .CK(clock), .Q(U72_DATA1_24), .QN(n34)
         );
  DFF_X1 temp_yVal_reg_25_ ( .D(n2656), .CK(clock), .Q(U72_DATA1_25), .QN(n33)
         );
  DFF_X1 temp_yVal_reg_26_ ( .D(n2657), .CK(clock), .Q(U72_DATA1_26), .QN(n32)
         );
  DFF_X1 temp_yVal_reg_27_ ( .D(n2658), .CK(clock), .Q(U72_DATA1_27), .QN(n31)
         );
  DFF_X1 temp_yVal_reg_28_ ( .D(n2659), .CK(clock), .Q(U72_DATA1_28), .QN(n30)
         );
  DFF_X1 op_yVal1_reg_47_ ( .D(U94_Z_47), .CK(clock), .Q(op_yVal1[47]) );
  DFF_X1 op_yVal1_reg_46_ ( .D(U94_Z_46), .CK(clock), .Q(op_yVal1[46]) );
  DFF_X1 op_yVal1_reg_45_ ( .D(U94_Z_45), .CK(clock), .Q(op_yVal1[45]) );
  DFF_X1 op_yVal1_reg_44_ ( .D(U94_Z_44), .CK(clock), .Q(op_yVal1[44]) );
  DFF_X1 op_yVal1_reg_43_ ( .D(U94_Z_43), .CK(clock), .Q(op_yVal1[43]) );
  DFF_X1 op_yVal1_reg_42_ ( .D(U94_Z_42), .CK(clock), .Q(op_yVal1[42]) );
  DFF_X1 op_yVal1_reg_41_ ( .D(U94_Z_41), .CK(clock), .Q(op_yVal1[41]) );
  DFF_X1 op_yVal1_reg_40_ ( .D(U94_Z_40), .CK(clock), .Q(op_yVal1[40]) );
  DFF_X1 op_yVal1_reg_39_ ( .D(U94_Z_39), .CK(clock), .Q(op_yVal1[39]) );
  DFF_X1 op_yVal1_reg_38_ ( .D(U94_Z_38), .CK(clock), .Q(op_yVal1[38]) );
  DFF_X1 op_yVal1_reg_37_ ( .D(U94_Z_37), .CK(clock), .Q(op_yVal1[37]) );
  DFF_X1 op_yVal1_reg_36_ ( .D(U94_Z_36), .CK(clock), .Q(op_yVal1[36]) );
  DFF_X1 op_yVal1_reg_35_ ( .D(U94_Z_35), .CK(clock), .Q(op_yVal1[35]) );
  DFF_X1 op_yVal1_reg_34_ ( .D(U94_Z_34), .CK(clock), .Q(op_yVal1[34]) );
  DFF_X1 op_yVal1_reg_33_ ( .D(U94_Z_33), .CK(clock), .Q(op_yVal1[33]) );
  DFF_X1 op_yVal1_reg_32_ ( .D(U94_Z_32), .CK(clock), .Q(op_yVal1[32]) );
  DFF_X1 op_yVal1_reg_31_ ( .D(U94_Z_31), .CK(clock), .Q(op_yVal1[31]) );
  DFF_X1 op_yVal1_reg_30_ ( .D(U94_Z_30), .CK(clock), .Q(op_yVal1[30]) );
  DFF_X1 op_yVal1_reg_29_ ( .D(U94_Z_29), .CK(clock), .Q(op_yVal1[29]) );
  DFF_X1 op_yVal1_reg_28_ ( .D(U94_Z_28), .CK(clock), .Q(op_yVal1[28]) );
  DFF_X1 op_yVal1_reg_27_ ( .D(U94_Z_27), .CK(clock), .Q(op_yVal1[27]) );
  DFF_X1 op_yVal1_reg_26_ ( .D(U94_Z_26), .CK(clock), .Q(op_yVal1[26]) );
  DFF_X1 op_yVal1_reg_25_ ( .D(U94_Z_25), .CK(clock), .Q(op_yVal1[25]) );
  DFF_X1 op_yVal1_reg_24_ ( .D(U94_Z_24), .CK(clock), .Q(op_yVal1[24]) );
  DFF_X1 op_yVal1_reg_23_ ( .D(U94_Z_23), .CK(clock), .Q(op_yVal1[23]) );
  DFF_X1 op_yVal1_reg_22_ ( .D(U94_Z_22), .CK(clock), .Q(op_yVal1[22]) );
  DFF_X1 op_yVal1_reg_21_ ( .D(U94_Z_21), .CK(clock), .Q(op_yVal1[21]) );
  DFF_X1 op_yVal1_reg_20_ ( .D(U94_Z_20), .CK(clock), .Q(op_yVal1[20]) );
  DFF_X1 op_yVal1_reg_19_ ( .D(U94_Z_19), .CK(clock), .Q(op_yVal1[19]) );
  DFF_X1 op_yVal1_reg_18_ ( .D(U94_Z_18), .CK(clock), .Q(op_yVal1[18]) );
  DFF_X1 op_yVal1_reg_17_ ( .D(U94_Z_17), .CK(clock), .Q(op_yVal1[17]) );
  DFF_X1 op_yVal1_reg_16_ ( .D(U94_Z_16), .CK(clock), .Q(op_yVal1[16]) );
  DFF_X1 op_yVal1_reg_15_ ( .D(U94_Z_15), .CK(clock), .Q(op_yVal1[15]) );
  DFF_X1 op_yVal1_reg_14_ ( .D(U94_Z_14), .CK(clock), .Q(op_yVal1[14]) );
  DFF_X1 op_yVal1_reg_13_ ( .D(U94_Z_13), .CK(clock), .Q(op_yVal1[13]) );
  DFF_X1 op_yVal1_reg_12_ ( .D(U94_Z_12), .CK(clock), .Q(op_yVal1[12]) );
  DFF_X1 op_yVal1_reg_11_ ( .D(U94_Z_11), .CK(clock), .Q(op_yVal1[11]) );
  DFF_X1 op_yVal1_reg_10_ ( .D(U94_Z_10), .CK(clock), .Q(op_yVal1[10]) );
  DFF_X1 op_yVal1_reg_9_ ( .D(U94_Z_9), .CK(clock), .Q(op_yVal1[9]) );
  DFF_X1 op_yVal1_reg_8_ ( .D(U94_Z_8), .CK(clock), .Q(op_yVal1[8]) );
  DFF_X1 op_yVal1_reg_7_ ( .D(U94_Z_7), .CK(clock), .Q(op_yVal1[7]) );
  DFF_X1 op_yVal1_reg_6_ ( .D(U94_Z_6), .CK(clock), .Q(op_yVal1[6]) );
  DFF_X1 op_yVal1_reg_5_ ( .D(U94_Z_5), .CK(clock), .Q(op_yVal1[5]) );
  DFF_X1 op_yVal1_reg_4_ ( .D(U94_Z_4), .CK(clock), .Q(op_yVal1[4]) );
  DFF_X1 op_yVal1_reg_3_ ( .D(U94_Z_3), .CK(clock), .Q(op_yVal1[3]) );
  DFF_X1 op_yVal1_reg_2_ ( .D(U94_Z_2), .CK(clock), .Q(op_yVal1[2]) );
  DFF_X1 op_yVal1_reg_1_ ( .D(U94_Z_1), .CK(clock), .Q(op_yVal1[1]) );
  DFF_X1 op_yVal1_reg_0_ ( .D(U94_Z_0), .CK(clock), .Q(op_yVal1[0]) );
  DFF_X1 op_yVal2_reg_47_ ( .D(U93_Z_47), .CK(clock), .Q(op_yVal2[47]) );
  DFF_X1 op_yVal2_reg_46_ ( .D(U93_Z_46), .CK(clock), .Q(op_yVal2[46]) );
  DFF_X1 op_yVal2_reg_45_ ( .D(U93_Z_45), .CK(clock), .Q(op_yVal2[45]) );
  DFF_X1 op_yVal2_reg_44_ ( .D(U93_Z_44), .CK(clock), .Q(op_yVal2[44]) );
  DFF_X1 op_yVal2_reg_43_ ( .D(U93_Z_43), .CK(clock), .Q(op_yVal2[43]) );
  DFF_X1 op_yVal2_reg_42_ ( .D(U93_Z_42), .CK(clock), .Q(op_yVal2[42]) );
  DFF_X1 op_yVal2_reg_41_ ( .D(U93_Z_41), .CK(clock), .Q(op_yVal2[41]) );
  DFF_X1 op_yVal2_reg_40_ ( .D(U93_Z_40), .CK(clock), .Q(op_yVal2[40]) );
  DFF_X1 op_yVal2_reg_39_ ( .D(U93_Z_39), .CK(clock), .Q(op_yVal2[39]) );
  DFF_X1 op_yVal2_reg_38_ ( .D(U93_Z_38), .CK(clock), .Q(op_yVal2[38]) );
  DFF_X1 op_yVal2_reg_37_ ( .D(U93_Z_37), .CK(clock), .Q(op_yVal2[37]) );
  DFF_X1 op_yVal2_reg_36_ ( .D(U93_Z_36), .CK(clock), .Q(op_yVal2[36]) );
  DFF_X1 op_yVal2_reg_35_ ( .D(U93_Z_35), .CK(clock), .Q(op_yVal2[35]) );
  DFF_X1 op_yVal2_reg_34_ ( .D(U93_Z_34), .CK(clock), .Q(op_yVal2[34]) );
  DFF_X1 op_yVal2_reg_33_ ( .D(U93_Z_33), .CK(clock), .Q(op_yVal2[33]) );
  DFF_X1 op_yVal2_reg_32_ ( .D(U93_Z_32), .CK(clock), .Q(op_yVal2[32]) );
  DFF_X1 op_yVal2_reg_31_ ( .D(U93_Z_31), .CK(clock), .Q(op_yVal2[31]) );
  DFF_X1 op_yVal2_reg_30_ ( .D(U93_Z_30), .CK(clock), .Q(op_yVal2[30]) );
  DFF_X1 op_yVal2_reg_29_ ( .D(U93_Z_29), .CK(clock), .Q(op_yVal2[29]) );
  DFF_X1 op_yVal2_reg_28_ ( .D(U93_Z_28), .CK(clock), .Q(op_yVal2[28]) );
  DFF_X1 op_yVal2_reg_27_ ( .D(U93_Z_27), .CK(clock), .Q(op_yVal2[27]) );
  DFF_X1 op_yVal2_reg_26_ ( .D(U93_Z_26), .CK(clock), .Q(op_yVal2[26]) );
  DFF_X1 op_yVal2_reg_25_ ( .D(U93_Z_25), .CK(clock), .Q(op_yVal2[25]) );
  DFF_X1 op_yVal2_reg_24_ ( .D(U93_Z_24), .CK(clock), .Q(op_yVal2[24]) );
  DFF_X1 op_yVal2_reg_23_ ( .D(U93_Z_23), .CK(clock), .Q(op_yVal2[23]) );
  DFF_X1 op_yVal2_reg_22_ ( .D(U93_Z_22), .CK(clock), .Q(op_yVal2[22]) );
  DFF_X1 op_yVal2_reg_21_ ( .D(U93_Z_21), .CK(clock), .Q(op_yVal2[21]) );
  DFF_X1 op_yVal2_reg_20_ ( .D(U93_Z_20), .CK(clock), .Q(op_yVal2[20]) );
  DFF_X1 op_yVal2_reg_19_ ( .D(U93_Z_19), .CK(clock), .Q(op_yVal2[19]) );
  DFF_X1 op_yVal2_reg_18_ ( .D(U93_Z_18), .CK(clock), .Q(op_yVal2[18]) );
  DFF_X1 op_yVal2_reg_17_ ( .D(U93_Z_17), .CK(clock), .Q(op_yVal2[17]) );
  DFF_X1 op_yVal2_reg_16_ ( .D(U93_Z_16), .CK(clock), .Q(op_yVal2[16]) );
  DFF_X1 op_yVal2_reg_15_ ( .D(U93_Z_15), .CK(clock), .Q(op_yVal2[15]) );
  DFF_X1 op_yVal2_reg_14_ ( .D(U93_Z_14), .CK(clock), .Q(op_yVal2[14]) );
  DFF_X1 op_yVal2_reg_13_ ( .D(U93_Z_13), .CK(clock), .Q(op_yVal2[13]) );
  DFF_X1 op_yVal2_reg_12_ ( .D(U93_Z_12), .CK(clock), .Q(op_yVal2[12]) );
  DFF_X1 op_yVal2_reg_11_ ( .D(U93_Z_11), .CK(clock), .Q(op_yVal2[11]) );
  DFF_X1 op_yVal2_reg_10_ ( .D(U93_Z_10), .CK(clock), .Q(op_yVal2[10]) );
  DFF_X1 op_yVal2_reg_9_ ( .D(U93_Z_9), .CK(clock), .Q(op_yVal2[9]) );
  DFF_X1 op_yVal2_reg_8_ ( .D(U93_Z_8), .CK(clock), .Q(op_yVal2[8]) );
  DFF_X1 op_yVal2_reg_7_ ( .D(U93_Z_7), .CK(clock), .Q(op_yVal2[7]) );
  DFF_X1 op_yVal2_reg_6_ ( .D(U93_Z_6), .CK(clock), .Q(op_yVal2[6]) );
  DFF_X1 op_yVal2_reg_5_ ( .D(U93_Z_5), .CK(clock), .Q(op_yVal2[5]) );
  DFF_X1 op_yVal2_reg_4_ ( .D(U93_Z_4), .CK(clock), .Q(op_yVal2[4]) );
  DFF_X1 op_yVal2_reg_3_ ( .D(U93_Z_3), .CK(clock), .Q(op_yVal2[3]) );
  DFF_X1 op_yVal2_reg_2_ ( .D(U93_Z_2), .CK(clock), .Q(op_yVal2[2]) );
  DFF_X1 op_yVal2_reg_1_ ( .D(U93_Z_1), .CK(clock), .Q(op_yVal2[1]) );
  DFF_X1 op_yVal2_reg_0_ ( .D(U93_Z_0), .CK(clock), .Q(op_yVal2[0]) );
  DFF_X1 op_EX_EN_reg ( .D(U92_Z_0), .CK(clock), .Q(op_EX_EN) );
  DFF_X1 op_y_row_reg_15_ ( .D(U91_Z_15), .CK(clock), .Q(op_y_row[15]) );
  DFF_X1 op_y_row_reg_14_ ( .D(U91_Z_14), .CK(clock), .Q(op_y_row[14]) );
  DFF_X1 op_y_row_reg_13_ ( .D(U91_Z_13), .CK(clock), .Q(op_y_row[13]) );
  DFF_X1 op_y_row_reg_12_ ( .D(U91_Z_12), .CK(clock), .Q(op_y_row[12]) );
  DFF_X1 op_y_row_reg_11_ ( .D(U91_Z_11), .CK(clock), .Q(op_y_row[11]) );
  DFF_X1 op_y_row_reg_10_ ( .D(U91_Z_10), .CK(clock), .Q(op_y_row[10]) );
  DFF_X1 op_y_row_reg_9_ ( .D(U91_Z_9), .CK(clock), .Q(op_y_row[9]) );
  DFF_X1 op_y_row_reg_8_ ( .D(U91_Z_8), .CK(clock), .Q(op_y_row[8]) );
  DFF_X1 op_y_row_reg_7_ ( .D(U91_Z_7), .CK(clock), .Q(op_y_row[7]) );
  DFF_X1 op_y_row_reg_6_ ( .D(U91_Z_6), .CK(clock), .Q(op_y_row[6]) );
  DFF_X1 op_y_row_reg_5_ ( .D(U91_Z_5), .CK(clock), .Q(op_y_row[5]) );
  DFF_X1 op_y_row_reg_4_ ( .D(U91_Z_4), .CK(clock), .Q(op_y_row[4]) );
  DFF_X1 op_y_row_reg_3_ ( .D(U91_Z_3), .CK(clock), .Q(op_y_row[3]) );
  DFF_X1 op_y_row_reg_2_ ( .D(U91_Z_2), .CK(clock), .Q(op_y_row[2]) );
  DFF_X1 op_y_row_reg_1_ ( .D(U91_Z_1), .CK(clock), .Q(op_y_row[1]) );
  DFF_X1 op_y_row_reg_0_ ( .D(U91_Z_0), .CK(clock), .Q(op_y_row[0]) );
  DFF_X1 op_DataEN_reg ( .D(U90_Z_0), .CK(clock), .Q(op_DataEN) );
  DFF_X1 op_yAddrDiag_reg_10_ ( .D(n60), .CK(clock), .Q(op_yAddrDiag[10]) );
  DFF_X1 op_yAddrDiag_reg_9_ ( .D(n61), .CK(clock), .Q(op_yAddrDiag[9]) );
  DFF_X1 op_yAddrDiag_reg_8_ ( .D(n62), .CK(clock), .Q(op_yAddrDiag[8]) );
  DFF_X1 op_yAddrDiag_reg_7_ ( .D(n63), .CK(clock), .Q(op_yAddrDiag[7]) );
  DFF_X1 op_yAddrDiag_reg_6_ ( .D(n64), .CK(clock), .Q(op_yAddrDiag[6]) );
  DFF_X1 op_yAddrDiag_reg_5_ ( .D(n65), .CK(clock), .Q(op_yAddrDiag[5]) );
  DFF_X1 op_yAddrDiag_reg_4_ ( .D(n66), .CK(clock), .Q(op_yAddrDiag[4]) );
  DFF_X1 op_yAddrDiag_reg_3_ ( .D(n67), .CK(clock), .Q(op_yAddrDiag[3]) );
  DFF_X1 op_yAddrDiag_reg_2_ ( .D(n68), .CK(clock), .Q(op_yAddrDiag[2]) );
  DFF_X1 op_yAddrDiag_reg_1_ ( .D(n69), .CK(clock), .Q(op_yAddrDiag[1]) );
  DFF_X1 op_yAddrDiag_reg_0_ ( .D(n70), .CK(clock), .Q(op_yAddrDiag[0]) );
  DFF_X1 op_yAddrNonDiag_reg_10_ ( .D(n2627), .CK(clock), .Q(
        op_yAddrNonDiag[10]) );
  DFF_X1 op_yAddrNonDiag_reg_9_ ( .D(n2626), .CK(clock), .Q(op_yAddrNonDiag[9]) );
  DFF_X1 op_yAddrNonDiag_reg_8_ ( .D(n2625), .CK(clock), .Q(op_yAddrNonDiag[8]) );
  DFF_X1 op_yAddrNonDiag_reg_7_ ( .D(n2624), .CK(clock), .Q(op_yAddrNonDiag[7]) );
  DFF_X1 op_yAddrNonDiag_reg_6_ ( .D(n2623), .CK(clock), .Q(op_yAddrNonDiag[6]) );
  DFF_X1 op_yAddrNonDiag_reg_5_ ( .D(n2622), .CK(clock), .Q(op_yAddrNonDiag[5]) );
  DFF_X1 op_yAddrNonDiag_reg_4_ ( .D(n2621), .CK(clock), .Q(op_yAddrNonDiag[4]) );
  DFF_X1 op_yAddrNonDiag_reg_3_ ( .D(n2620), .CK(clock), .Q(op_yAddrNonDiag[3]) );
  DFF_X1 op_yAddrNonDiag_reg_2_ ( .D(n2619), .CK(clock), .Q(op_yAddrNonDiag[2]) );
  DFF_X1 op_yAddrNonDiag_reg_1_ ( .D(n2618), .CK(clock), .Q(op_yAddrNonDiag[1]) );
  DFF_X1 op_yAddrNonDiag_reg_0_ ( .D(n2617), .CK(clock), .Q(op_yAddrNonDiag[0]) );
  DFF_X2 op_oneHotDiag_reg_3_ ( .D(n2616), .CK(clock), .Q(op_oneHotDiag[3]), 
        .QN(n153) );
  DFF_X2 op_oneHotDiag_reg_2_ ( .D(n2615), .CK(clock), .Q(op_oneHotDiag[2]), 
        .QN(n154) );
  DFF_X1 op_oneHotDiag_reg_1_ ( .D(n2614), .CK(clock), .Q(op_oneHotDiag[1]) );
  DFF_X1 op_oneHotDiag_reg_0_ ( .D(n71), .CK(clock), .Q(op_oneHotDiag[0]) );
  NAND2_X2 U5 ( .A1(op_oneHotDiag[1]), .A2(n72), .ZN(n630) );
  OAI22_X2 U6 ( .A1(n632), .A2(n154), .B1(n3281), .B2(n629), .ZN(n2615) );
  OAI22_X2 U7 ( .A1(n632), .A2(n153), .B1(n3216), .B2(n629), .ZN(n2616) );
  NAND2_X2 U8 ( .A1(n632), .A2(reset), .ZN(n629) );
  AOI221_X2 U10 ( .B1(n3291), .B2(n85), .C1(op_yAddrNonDiag[0]), .C2(n7), .A(
        n637), .ZN(n636) );
  AOI221_X2 U11 ( .B1(n639), .B2(yAddrIn2[0]), .C1(n640), .C2(yAddrIn1[0]), 
        .A(n641), .ZN(n638) );
  AOI221_X2 U13 ( .B1(yAddrIn2[0]), .B2(n644), .C1(yAddrIn1[0]), .C2(n645), 
        .A(n646), .ZN(n633) );
  AOI221_X2 U15 ( .B1(n3291), .B2(n84), .C1(op_yAddrNonDiag[1]), .C2(n7), .A(
        n637), .ZN(n649) );
  AOI221_X2 U16 ( .B1(n639), .B2(yAddrIn2[1]), .C1(n640), .C2(yAddrIn1[1]), 
        .A(n641), .ZN(n650) );
  AOI221_X2 U18 ( .B1(yAddrIn2[1]), .B2(n644), .C1(yAddrIn1[1]), .C2(n645), 
        .A(n646), .ZN(n647) );
  AOI221_X2 U20 ( .B1(n3291), .B2(n83), .C1(op_yAddrNonDiag[2]), .C2(n7), .A(
        n637), .ZN(n653) );
  AOI221_X2 U21 ( .B1(n639), .B2(yAddrIn2[2]), .C1(n640), .C2(yAddrIn1[2]), 
        .A(n641), .ZN(n654) );
  AOI221_X2 U23 ( .B1(yAddrIn2[2]), .B2(n644), .C1(yAddrIn1[2]), .C2(n645), 
        .A(n646), .ZN(n651) );
  AOI221_X2 U25 ( .B1(n3291), .B2(n82), .C1(op_yAddrNonDiag[3]), .C2(n7), .A(
        n637), .ZN(n657) );
  AOI221_X2 U26 ( .B1(n639), .B2(yAddrIn2[3]), .C1(n640), .C2(yAddrIn1[3]), 
        .A(n641), .ZN(n658) );
  AOI221_X2 U28 ( .B1(yAddrIn2[3]), .B2(n644), .C1(yAddrIn1[3]), .C2(n645), 
        .A(n646), .ZN(n655) );
  AOI221_X2 U30 ( .B1(n3291), .B2(n81), .C1(op_yAddrNonDiag[4]), .C2(n7), .A(
        n637), .ZN(n661) );
  AOI221_X2 U31 ( .B1(n639), .B2(yAddrIn2[4]), .C1(n640), .C2(yAddrIn1[4]), 
        .A(n641), .ZN(n662) );
  AOI221_X2 U33 ( .B1(yAddrIn2[4]), .B2(n644), .C1(yAddrIn1[4]), .C2(n645), 
        .A(n646), .ZN(n659) );
  AOI221_X2 U35 ( .B1(n3291), .B2(n80), .C1(op_yAddrNonDiag[5]), .C2(n7), .A(
        n637), .ZN(n665) );
  AOI221_X2 U36 ( .B1(n639), .B2(yAddrIn2[5]), .C1(n640), .C2(yAddrIn1[5]), 
        .A(n641), .ZN(n666) );
  AOI221_X2 U38 ( .B1(yAddrIn2[5]), .B2(n644), .C1(yAddrIn1[5]), .C2(n645), 
        .A(n646), .ZN(n663) );
  AOI221_X2 U40 ( .B1(n3291), .B2(n79), .C1(op_yAddrNonDiag[6]), .C2(n7), .A(
        n637), .ZN(n669) );
  AOI221_X2 U41 ( .B1(n639), .B2(yAddrIn2[6]), .C1(n640), .C2(yAddrIn1[6]), 
        .A(n641), .ZN(n670) );
  AOI221_X2 U43 ( .B1(yAddrIn2[6]), .B2(n644), .C1(yAddrIn1[6]), .C2(n645), 
        .A(n646), .ZN(n667) );
  AOI221_X2 U45 ( .B1(n3291), .B2(n78), .C1(op_yAddrNonDiag[7]), .C2(n7), .A(
        n637), .ZN(n673) );
  AOI221_X2 U46 ( .B1(n639), .B2(yAddrIn2[7]), .C1(n640), .C2(yAddrIn1[7]), 
        .A(n641), .ZN(n674) );
  AOI221_X2 U48 ( .B1(yAddrIn2[7]), .B2(n644), .C1(yAddrIn1[7]), .C2(n645), 
        .A(n646), .ZN(n671) );
  AOI221_X2 U50 ( .B1(n3291), .B2(n77), .C1(op_yAddrNonDiag[8]), .C2(n7), .A(
        n637), .ZN(n677) );
  AOI221_X2 U51 ( .B1(n639), .B2(yAddrIn2[8]), .C1(n640), .C2(yAddrIn1[8]), 
        .A(n641), .ZN(n678) );
  AOI221_X2 U53 ( .B1(yAddrIn2[8]), .B2(n644), .C1(yAddrIn1[8]), .C2(n645), 
        .A(n646), .ZN(n675) );
  AOI221_X2 U55 ( .B1(n3291), .B2(n76), .C1(op_yAddrNonDiag[9]), .C2(n7), .A(
        n637), .ZN(n681) );
  AOI221_X2 U56 ( .B1(n639), .B2(yAddrIn2[9]), .C1(n640), .C2(yAddrIn1[9]), 
        .A(n641), .ZN(n682) );
  AOI221_X2 U58 ( .B1(yAddrIn2[9]), .B2(n644), .C1(yAddrIn1[9]), .C2(n645), 
        .A(n646), .ZN(n679) );
  AOI221_X2 U60 ( .B1(n3291), .B2(n75), .C1(op_yAddrNonDiag[10]), .C2(n7), .A(
        n637), .ZN(n685) );
  AOI221_X2 U62 ( .B1(n639), .B2(yAddrIn2[10]), .C1(n640), .C2(yAddrIn1[10]), 
        .A(n641), .ZN(n686) );
  AOI221_X2 U64 ( .B1(n690), .B2(n136), .C1(n88), .C2(n122), .A(n691), .ZN(
        n689) );
  NOR3_X2 U65 ( .A1(n692), .A2(n693), .A3(n137), .ZN(n691) );
  NOR3_X2 U67 ( .A1(n111), .A2(n112), .A3(n699), .ZN(n694) );
  NAND3_X2 U68 ( .A1(n700), .A2(n701), .A3(n702), .ZN(n639) );
  NAND4_X2 U70 ( .A1(n93), .A2(n706), .A3(n101), .A4(n707), .ZN(n705) );
  NAND4_X2 U71 ( .A1(n708), .A2(n709), .A3(n710), .A4(n711), .ZN(n703) );
  NOR4_X2 U75 ( .A1(n718), .A2(n719), .A3(n720), .A4(n721), .ZN(n716) );
  NOR2_X2 U76 ( .A1(n722), .A2(n723), .ZN(n721) );
  AOI221_X2 U80 ( .B1(yAddrIn2[10]), .B2(n644), .C1(yAddrIn1[10]), .C2(n645), 
        .A(n646), .ZN(n683) );
  AOI221_X2 U82 ( .B1(n87), .B2(n115), .C1(n89), .C2(n120), .A(n731), .ZN(n730) );
  NOR3_X2 U83 ( .A1(n692), .A2(n116), .A3(n732), .ZN(n731) );
  NOR3_X2 U85 ( .A1(n111), .A2(n105), .A3(n736), .ZN(n733) );
  NOR2_X2 U86 ( .A1(n132), .A2(n737), .ZN(n696) );
  NAND3_X2 U87 ( .A1(n738), .A2(n739), .A3(n740), .ZN(n644) );
  NAND4_X2 U89 ( .A1(n743), .A2(n744), .A3(n101), .A4(n707), .ZN(n742) );
  NAND4_X2 U90 ( .A1(n746), .A2(n98), .A3(n747), .A4(n748), .ZN(n741) );
  AOI221_X2 U92 ( .B1(n72), .B2(op_yAddrDiag[0]), .C1(n632), .C2(yAddrIn1[0]), 
        .A(n3300), .ZN(n753) );
  AOI221_X2 U93 ( .B1(n72), .B2(op_yAddrDiag[1]), .C1(n632), .C2(yAddrIn1[1]), 
        .A(n3300), .ZN(n754) );
  AOI221_X2 U94 ( .B1(n72), .B2(op_yAddrDiag[2]), .C1(n632), .C2(yAddrIn1[2]), 
        .A(n3300), .ZN(n755) );
  AOI221_X2 U95 ( .B1(n72), .B2(op_yAddrDiag[3]), .C1(n632), .C2(yAddrIn1[3]), 
        .A(n3300), .ZN(n756) );
  AOI221_X2 U96 ( .B1(n72), .B2(op_yAddrDiag[4]), .C1(n632), .C2(yAddrIn1[4]), 
        .A(n3300), .ZN(n757) );
  AOI221_X2 U97 ( .B1(n72), .B2(op_yAddrDiag[5]), .C1(n632), .C2(yAddrIn1[5]), 
        .A(n3300), .ZN(n758) );
  AOI221_X2 U98 ( .B1(n72), .B2(op_yAddrDiag[6]), .C1(n632), .C2(yAddrIn1[6]), 
        .A(n3300), .ZN(n759) );
  AOI221_X2 U99 ( .B1(n72), .B2(op_yAddrDiag[7]), .C1(n632), .C2(yAddrIn1[7]), 
        .A(n3300), .ZN(n760) );
  AOI221_X2 U100 ( .B1(n72), .B2(op_yAddrDiag[8]), .C1(n632), .C2(yAddrIn1[8]), 
        .A(n3300), .ZN(n761) );
  AOI221_X2 U101 ( .B1(n72), .B2(op_yAddrDiag[9]), .C1(n632), .C2(yAddrIn1[9]), 
        .A(n3300), .ZN(n762) );
  AOI221_X2 U102 ( .B1(n72), .B2(op_yAddrDiag[10]), .C1(n632), .C2(
        yAddrIn1[10]), .A(n3300), .ZN(n763) );
  NAND4_X2 U105 ( .A1(n768), .A2(n769), .A3(n770), .A4(n771), .ZN(n767) );
  NOR3_X2 U106 ( .A1(n772), .A2(n773), .A3(n774), .ZN(n771) );
  NOR2_X2 U110 ( .A1(n780), .A2(n5), .ZN(n779) );
  NOR2_X2 U112 ( .A1(n3303), .A2(n722), .ZN(n720) );
  NAND2_X2 U116 ( .A1(op_oneHotNonDiag[1]), .A2(n7), .ZN(n787) );
  NOR4_X2 U117 ( .A1(n788), .A2(n10), .A3(n789), .A4(n790), .ZN(n785) );
  NOR2_X2 U121 ( .A1(n3305), .A2(n722), .ZN(n719) );
  OAI221_X2 U122 ( .B1(n801), .B2(n3286), .C1(n777), .C2(n3307), .A(n803), 
        .ZN(n788) );
  NOR2_X2 U124 ( .A1(n804), .A2(n805), .ZN(n801) );
  NAND2_X2 U126 ( .A1(op_oneHotNonDiag[2]), .A2(n7), .ZN(n807) );
  NOR4_X2 U127 ( .A1(n808), .A2(n809), .A3(n810), .A4(n6), .ZN(n806) );
  OAI22_X2 U130 ( .A1(n3290), .A2(n102), .B1(n777), .B2(n815), .ZN(n809) );
  OAI221_X2 U131 ( .B1(n775), .B2(n747), .C1(n710), .C2(n776), .A(n816), .ZN(
        n808) );
  NAND2_X2 U133 ( .A1(n818), .A2(n819), .ZN(n2630) );
  NAND2_X2 U135 ( .A1(n822), .A2(reset), .ZN(n786) );
  OAI221_X2 U136 ( .B1(n711), .B2(n776), .C1(n3286), .C2(n823), .A(n824), .ZN(
        n821) );
  OAI221_X2 U138 ( .B1(n3290), .B2(n825), .C1(n3281), .C2(n707), .A(n826), 
        .ZN(n820) );
  NAND2_X2 U140 ( .A1(n793), .A2(n777), .ZN(n827) );
  NAND2_X2 U141 ( .A1(n9), .A2(n130), .ZN(n777) );
  NAND2_X2 U142 ( .A1(op_oneHotNonDiag[3]), .A2(n7), .ZN(n818) );
  OAI221_X2 U145 ( .B1(n832), .B2(n3274), .C1(n3309), .C2(n58), .A(n835), .ZN(
        n2631) );
  AOI221_X2 U148 ( .B1(ymem_data2[128]), .B2(n3276), .C1(ymem_data2[192]), 
        .C2(n3297), .A(n843), .ZN(n841) );
  OAI22_X2 U149 ( .A1(n3305), .A2(n562), .B1(n3303), .B2(n626), .ZN(n843) );
  AOI221_X2 U150 ( .B1(ymem_data1[128]), .B2(n3292), .C1(ymem_data1[192]), 
        .C2(n3257), .A(n844), .ZN(n840) );
  OAI22_X2 U151 ( .A1(n3307), .A2(n370), .B1(n778), .B2(n434), .ZN(n844) );
  AOI221_X2 U153 ( .B1(ymem_data2[128]), .B2(n3270), .C1(ymem_data2[192]), 
        .C2(n3268), .A(n850), .ZN(n846) );
  OAI22_X2 U154 ( .A1(n3266), .A2(n562), .B1(n3264), .B2(n626), .ZN(n850) );
  AOI221_X2 U155 ( .B1(ymem_data1[0]), .B2(n3263), .C1(ymem_data1[64]), .C2(
        n3261), .A(n855), .ZN(n845) );
  AOI221_X2 U158 ( .B1(ymem_data1[0]), .B2(n3293), .C1(ymem_data2[192]), .C2(
        n3253), .A(n861), .ZN(n859) );
  OAI22_X2 U159 ( .A1(n3251), .A2(n370), .B1(n306), .B2(n3249), .ZN(n861) );
  OAI22_X2 U162 ( .A1(n3240), .A2(n562), .B1(n99), .B2(n498), .ZN(n868) );
  OAI221_X2 U165 ( .B1(n872), .B2(n3275), .C1(n3309), .C2(n57), .A(n873), .ZN(
        n2632) );
  AOI221_X2 U168 ( .B1(ymem_data2[129]), .B2(n3276), .C1(ymem_data2[193]), 
        .C2(n3297), .A(n879), .ZN(n878) );
  OAI22_X2 U169 ( .A1(n3305), .A2(n561), .B1(n3303), .B2(n625), .ZN(n879) );
  AOI221_X2 U170 ( .B1(ymem_data1[129]), .B2(n3292), .C1(ymem_data1[193]), 
        .C2(n3257), .A(n880), .ZN(n877) );
  OAI22_X2 U171 ( .A1(n3307), .A2(n369), .B1(n778), .B2(n433), .ZN(n880) );
  AOI221_X2 U173 ( .B1(ymem_data2[129]), .B2(n3270), .C1(ymem_data2[193]), 
        .C2(n3268), .A(n883), .ZN(n882) );
  OAI22_X2 U174 ( .A1(n3266), .A2(n561), .B1(n3264), .B2(n625), .ZN(n883) );
  AOI221_X2 U175 ( .B1(ymem_data1[1]), .B2(n3263), .C1(ymem_data1[65]), .C2(
        n3261), .A(n884), .ZN(n881) );
  OAI22_X2 U176 ( .A1(n3259), .A2(n241), .B1(n3255), .B2(n305), .ZN(n884) );
  AOI221_X2 U178 ( .B1(ymem_data1[1]), .B2(n3293), .C1(ymem_data2[193]), .C2(
        n3253), .A(n887), .ZN(n886) );
  OAI22_X2 U179 ( .A1(n862), .A2(n369), .B1(n3249), .B2(n305), .ZN(n887) );
  OAI22_X2 U182 ( .A1(n3240), .A2(n561), .B1(n99), .B2(n497), .ZN(n889) );
  OAI221_X2 U183 ( .B1(n3248), .B2(n305), .C1(n870), .C2(n369), .A(n890), .ZN(
        n888) );
  OAI221_X2 U185 ( .B1(n891), .B2(n3275), .C1(n3309), .C2(n56), .A(n892), .ZN(
        n2633) );
  AOI221_X2 U188 ( .B1(ymem_data2[130]), .B2(n3276), .C1(ymem_data2[194]), 
        .C2(n3297), .A(n898), .ZN(n897) );
  OAI22_X2 U189 ( .A1(n3305), .A2(n560), .B1(n3303), .B2(n624), .ZN(n898) );
  AOI221_X2 U190 ( .B1(ymem_data1[130]), .B2(n3292), .C1(ymem_data1[194]), 
        .C2(n3257), .A(n899), .ZN(n896) );
  OAI22_X2 U191 ( .A1(n3307), .A2(n368), .B1(n778), .B2(n432), .ZN(n899) );
  AOI221_X2 U193 ( .B1(ymem_data2[130]), .B2(n3270), .C1(ymem_data2[194]), 
        .C2(n3268), .A(n902), .ZN(n901) );
  OAI22_X2 U194 ( .A1(n3266), .A2(n560), .B1(n3264), .B2(n624), .ZN(n902) );
  AOI221_X2 U195 ( .B1(ymem_data1[2]), .B2(n3262), .C1(ymem_data1[66]), .C2(
        n3261), .A(n903), .ZN(n900) );
  OAI22_X2 U196 ( .A1(n3259), .A2(n240), .B1(n857), .B2(n304), .ZN(n903) );
  AOI221_X2 U198 ( .B1(ymem_data1[2]), .B2(n3293), .C1(ymem_data2[194]), .C2(
        n3253), .A(n906), .ZN(n905) );
  OAI22_X2 U199 ( .A1(n862), .A2(n368), .B1(n3249), .B2(n304), .ZN(n906) );
  OAI22_X2 U202 ( .A1(n869), .A2(n560), .B1(n99), .B2(n496), .ZN(n908) );
  OAI221_X2 U203 ( .B1(n3248), .B2(n304), .C1(n870), .C2(n368), .A(n909), .ZN(
        n907) );
  OAI221_X2 U205 ( .B1(n910), .B2(n3274), .C1(n3309), .C2(n55), .A(n911), .ZN(
        n2634) );
  AOI221_X2 U208 ( .B1(ymem_data2[131]), .B2(n3276), .C1(ymem_data2[195]), 
        .C2(n3297), .A(n917), .ZN(n916) );
  OAI22_X2 U209 ( .A1(n3305), .A2(n559), .B1(n3303), .B2(n623), .ZN(n917) );
  AOI221_X2 U210 ( .B1(ymem_data1[131]), .B2(n3292), .C1(ymem_data1[195]), 
        .C2(n3258), .A(n918), .ZN(n915) );
  OAI22_X2 U211 ( .A1(n3307), .A2(n367), .B1(n778), .B2(n431), .ZN(n918) );
  AOI221_X2 U213 ( .B1(ymem_data2[131]), .B2(n3270), .C1(ymem_data2[195]), 
        .C2(n3268), .A(n921), .ZN(n920) );
  OAI22_X2 U214 ( .A1(n3266), .A2(n559), .B1(n3264), .B2(n623), .ZN(n921) );
  AOI221_X2 U215 ( .B1(ymem_data1[3]), .B2(n3263), .C1(ymem_data1[67]), .C2(
        n3261), .A(n922), .ZN(n919) );
  OAI22_X2 U216 ( .A1(n3259), .A2(n239), .B1(n3255), .B2(n303), .ZN(n922) );
  AOI221_X2 U218 ( .B1(ymem_data1[3]), .B2(n3293), .C1(ymem_data2[195]), .C2(
        n860), .A(n925), .ZN(n924) );
  OAI22_X2 U219 ( .A1(n862), .A2(n367), .B1(n3248), .B2(n303), .ZN(n925) );
  OAI22_X2 U222 ( .A1(n869), .A2(n559), .B1(n99), .B2(n495), .ZN(n927) );
  OAI221_X2 U223 ( .B1(n3248), .B2(n303), .C1(n870), .C2(n367), .A(n928), .ZN(
        n926) );
  OAI221_X2 U225 ( .B1(n929), .B2(n3275), .C1(n3309), .C2(n54), .A(n930), .ZN(
        n2635) );
  AOI221_X2 U228 ( .B1(ymem_data2[132]), .B2(n3276), .C1(ymem_data2[196]), 
        .C2(n3297), .A(n936), .ZN(n935) );
  OAI22_X2 U229 ( .A1(n3305), .A2(n558), .B1(n3303), .B2(n622), .ZN(n936) );
  AOI221_X2 U230 ( .B1(ymem_data1[132]), .B2(n3292), .C1(ymem_data1[196]), 
        .C2(n3258), .A(n937), .ZN(n934) );
  OAI22_X2 U231 ( .A1(n3307), .A2(n366), .B1(n778), .B2(n430), .ZN(n937) );
  AOI221_X2 U233 ( .B1(ymem_data2[132]), .B2(n3270), .C1(ymem_data2[196]), 
        .C2(n3268), .A(n940), .ZN(n939) );
  OAI22_X2 U234 ( .A1(n3266), .A2(n558), .B1(n3264), .B2(n622), .ZN(n940) );
  AOI221_X2 U235 ( .B1(ymem_data1[4]), .B2(n3262), .C1(ymem_data1[68]), .C2(
        n3261), .A(n941), .ZN(n938) );
  OAI22_X2 U236 ( .A1(n3259), .A2(n238), .B1(n3255), .B2(n302), .ZN(n941) );
  AOI221_X2 U238 ( .B1(ymem_data1[4]), .B2(n3294), .C1(ymem_data2[196]), .C2(
        n860), .A(n944), .ZN(n943) );
  OAI22_X2 U242 ( .A1(n3240), .A2(n558), .B1(n99), .B2(n494), .ZN(n946) );
  OAI221_X2 U243 ( .B1(n3248), .B2(n302), .C1(n870), .C2(n366), .A(n947), .ZN(
        n945) );
  OAI221_X2 U245 ( .B1(n948), .B2(n3274), .C1(n3309), .C2(n53), .A(n949), .ZN(
        n2636) );
  AOI221_X2 U248 ( .B1(ymem_data2[133]), .B2(n3276), .C1(ymem_data2[197]), 
        .C2(n3297), .A(n955), .ZN(n954) );
  OAI22_X2 U249 ( .A1(n3305), .A2(n557), .B1(n3303), .B2(n621), .ZN(n955) );
  AOI221_X2 U250 ( .B1(ymem_data1[133]), .B2(n3292), .C1(ymem_data1[197]), 
        .C2(n3258), .A(n956), .ZN(n953) );
  OAI22_X2 U251 ( .A1(n3307), .A2(n365), .B1(n778), .B2(n429), .ZN(n956) );
  AOI221_X2 U253 ( .B1(ymem_data2[133]), .B2(n3270), .C1(ymem_data2[197]), 
        .C2(n3268), .A(n959), .ZN(n958) );
  OAI22_X2 U254 ( .A1(n3266), .A2(n557), .B1(n3264), .B2(n621), .ZN(n959) );
  AOI221_X2 U255 ( .B1(ymem_data1[5]), .B2(n3263), .C1(ymem_data1[69]), .C2(
        n3261), .A(n960), .ZN(n957) );
  OAI22_X2 U256 ( .A1(n856), .A2(n237), .B1(n3255), .B2(n301), .ZN(n960) );
  AOI221_X2 U258 ( .B1(ymem_data1[5]), .B2(n3293), .C1(ymem_data2[197]), .C2(
        n3253), .A(n963), .ZN(n962) );
  OAI22_X2 U259 ( .A1(n3251), .A2(n365), .B1(n863), .B2(n301), .ZN(n963) );
  OAI22_X2 U262 ( .A1(n869), .A2(n557), .B1(n99), .B2(n493), .ZN(n965) );
  OAI221_X2 U263 ( .B1(n863), .B2(n301), .C1(n870), .C2(n365), .A(n966), .ZN(
        n964) );
  OAI221_X2 U265 ( .B1(n967), .B2(n3274), .C1(n3309), .C2(n52), .A(n968), .ZN(
        n2637) );
  AOI221_X2 U268 ( .B1(ymem_data2[134]), .B2(n3276), .C1(ymem_data2[198]), 
        .C2(n3297), .A(n974), .ZN(n973) );
  OAI22_X2 U269 ( .A1(n3305), .A2(n556), .B1(n3303), .B2(n620), .ZN(n974) );
  AOI221_X2 U270 ( .B1(ymem_data1[134]), .B2(n3292), .C1(ymem_data1[198]), 
        .C2(n3258), .A(n975), .ZN(n972) );
  OAI22_X2 U271 ( .A1(n3307), .A2(n364), .B1(n778), .B2(n428), .ZN(n975) );
  AOI221_X2 U273 ( .B1(ymem_data2[134]), .B2(n3270), .C1(ymem_data2[198]), 
        .C2(n3268), .A(n978), .ZN(n977) );
  OAI22_X2 U274 ( .A1(n3266), .A2(n556), .B1(n3264), .B2(n620), .ZN(n978) );
  AOI221_X2 U275 ( .B1(ymem_data1[6]), .B2(n3262), .C1(ymem_data1[70]), .C2(
        n3261), .A(n979), .ZN(n976) );
  AOI221_X2 U278 ( .B1(ymem_data1[6]), .B2(n3294), .C1(ymem_data2[198]), .C2(
        n3253), .A(n982), .ZN(n981) );
  OAI22_X2 U279 ( .A1(n3251), .A2(n364), .B1(n863), .B2(n300), .ZN(n982) );
  OAI22_X2 U282 ( .A1(n869), .A2(n556), .B1(n99), .B2(n492), .ZN(n984) );
  OAI221_X2 U283 ( .B1(n863), .B2(n300), .C1(n870), .C2(n364), .A(n985), .ZN(
        n983) );
  OAI221_X2 U285 ( .B1(n986), .B2(n3275), .C1(n3309), .C2(n51), .A(n987), .ZN(
        n2638) );
  AOI221_X2 U288 ( .B1(ymem_data2[135]), .B2(n3276), .C1(ymem_data2[199]), 
        .C2(n3297), .A(n993), .ZN(n992) );
  OAI22_X2 U289 ( .A1(n3305), .A2(n555), .B1(n3303), .B2(n619), .ZN(n993) );
  AOI221_X2 U290 ( .B1(ymem_data1[135]), .B2(n3292), .C1(ymem_data1[199]), 
        .C2(n3258), .A(n994), .ZN(n991) );
  OAI22_X2 U291 ( .A1(n3307), .A2(n363), .B1(n778), .B2(n427), .ZN(n994) );
  OAI22_X2 U294 ( .A1(n3266), .A2(n555), .B1(n3264), .B2(n619), .ZN(n997) );
  AOI221_X2 U295 ( .B1(ymem_data1[7]), .B2(n3263), .C1(ymem_data1[71]), .C2(
        n3261), .A(n998), .ZN(n995) );
  OAI22_X2 U296 ( .A1(n856), .A2(n235), .B1(n3255), .B2(n299), .ZN(n998) );
  AOI221_X2 U298 ( .B1(ymem_data1[7]), .B2(n3294), .C1(ymem_data2[199]), .C2(
        n860), .A(n1001), .ZN(n1000) );
  OAI22_X2 U299 ( .A1(n862), .A2(n363), .B1(n863), .B2(n299), .ZN(n1001) );
  OAI22_X2 U302 ( .A1(n3240), .A2(n555), .B1(n99), .B2(n491), .ZN(n1003) );
  OAI221_X2 U303 ( .B1(n863), .B2(n299), .C1(n870), .C2(n363), .A(n1004), .ZN(
        n1002) );
  OAI221_X2 U305 ( .B1(n1005), .B2(n3275), .C1(n3309), .C2(n50), .A(n1006), 
        .ZN(n2639) );
  AOI221_X2 U308 ( .B1(ymem_data2[136]), .B2(n3276), .C1(ymem_data2[200]), 
        .C2(n3297), .A(n1012), .ZN(n1011) );
  OAI22_X2 U309 ( .A1(n3305), .A2(n554), .B1(n3303), .B2(n618), .ZN(n1012) );
  AOI221_X2 U310 ( .B1(ymem_data1[136]), .B2(n3292), .C1(ymem_data1[200]), 
        .C2(n3258), .A(n1013), .ZN(n1010) );
  OAI22_X2 U311 ( .A1(n3307), .A2(n362), .B1(n3284), .B2(n426), .ZN(n1013) );
  AOI221_X2 U313 ( .B1(ymem_data2[136]), .B2(n3270), .C1(ymem_data2[200]), 
        .C2(n3268), .A(n1016), .ZN(n1015) );
  OAI22_X2 U314 ( .A1(n3266), .A2(n554), .B1(n3264), .B2(n618), .ZN(n1016) );
  AOI221_X2 U315 ( .B1(ymem_data1[8]), .B2(n3262), .C1(ymem_data1[72]), .C2(
        n3261), .A(n1017), .ZN(n1014) );
  AOI221_X2 U318 ( .B1(ymem_data1[8]), .B2(n3293), .C1(ymem_data2[200]), .C2(
        n860), .A(n1020), .ZN(n1019) );
  OAI22_X2 U319 ( .A1(n3251), .A2(n362), .B1(n3248), .B2(n298), .ZN(n1020) );
  OAI22_X2 U322 ( .A1(n869), .A2(n554), .B1(n99), .B2(n490), .ZN(n1022) );
  OAI221_X2 U323 ( .B1(n863), .B2(n298), .C1(n3238), .C2(n362), .A(n1023), 
        .ZN(n1021) );
  OAI221_X2 U325 ( .B1(n1024), .B2(n3274), .C1(n3309), .C2(n49), .A(n1025), 
        .ZN(n2640) );
  AOI221_X2 U328 ( .B1(ymem_data2[137]), .B2(n3277), .C1(ymem_data2[201]), 
        .C2(n3296), .A(n1031), .ZN(n1030) );
  OAI22_X2 U329 ( .A1(n3305), .A2(n553), .B1(n3303), .B2(n617), .ZN(n1031) );
  AOI221_X2 U330 ( .B1(ymem_data1[137]), .B2(n3292), .C1(ymem_data1[201]), 
        .C2(n3258), .A(n1032), .ZN(n1029) );
  OAI22_X2 U331 ( .A1(n3307), .A2(n361), .B1(n3284), .B2(n425), .ZN(n1032) );
  AOI221_X2 U333 ( .B1(ymem_data2[137]), .B2(n3271), .C1(ymem_data2[201]), 
        .C2(n3268), .A(n1035), .ZN(n1034) );
  OAI22_X2 U334 ( .A1(n3266), .A2(n553), .B1(n3264), .B2(n617), .ZN(n1035) );
  AOI221_X2 U335 ( .B1(ymem_data1[9]), .B2(n3263), .C1(ymem_data1[73]), .C2(
        n3261), .A(n1036), .ZN(n1033) );
  OAI22_X2 U336 ( .A1(n856), .A2(n233), .B1(n3255), .B2(n297), .ZN(n1036) );
  AOI221_X2 U338 ( .B1(ymem_data1[9]), .B2(n3293), .C1(ymem_data2[201]), .C2(
        n860), .A(n1039), .ZN(n1038) );
  OAI22_X2 U339 ( .A1(n3251), .A2(n361), .B1(n863), .B2(n297), .ZN(n1039) );
  OAI22_X2 U342 ( .A1(n3240), .A2(n553), .B1(n99), .B2(n489), .ZN(n1041) );
  OAI221_X2 U343 ( .B1(n3248), .B2(n297), .C1(n870), .C2(n361), .A(n1042), 
        .ZN(n1040) );
  OAI221_X2 U345 ( .B1(n1043), .B2(n3275), .C1(n3309), .C2(n48), .A(n1044), 
        .ZN(n2641) );
  AOI221_X2 U348 ( .B1(ymem_data2[138]), .B2(n3277), .C1(ymem_data2[202]), 
        .C2(n3296), .A(n1050), .ZN(n1049) );
  OAI22_X2 U349 ( .A1(n3305), .A2(n552), .B1(n3303), .B2(n616), .ZN(n1050) );
  AOI221_X2 U350 ( .B1(ymem_data1[138]), .B2(n3292), .C1(ymem_data1[202]), 
        .C2(n3258), .A(n1051), .ZN(n1048) );
  OAI22_X2 U351 ( .A1(n3307), .A2(n360), .B1(n3284), .B2(n424), .ZN(n1051) );
  OAI22_X2 U354 ( .A1(n3266), .A2(n552), .B1(n3264), .B2(n616), .ZN(n1054) );
  AOI221_X2 U355 ( .B1(ymem_data1[10]), .B2(n3262), .C1(ymem_data1[74]), .C2(
        n854), .A(n1055), .ZN(n1052) );
  OAI22_X2 U356 ( .A1(n856), .A2(n232), .B1(n3255), .B2(n296), .ZN(n1055) );
  AOI221_X2 U358 ( .B1(ymem_data1[10]), .B2(n3294), .C1(ymem_data2[202]), .C2(
        n860), .A(n1058), .ZN(n1057) );
  OAI22_X2 U359 ( .A1(n3251), .A2(n360), .B1(n3248), .B2(n296), .ZN(n1058) );
  OAI22_X2 U362 ( .A1(n869), .A2(n552), .B1(n99), .B2(n488), .ZN(n1060) );
  OAI221_X2 U363 ( .B1(n3248), .B2(n296), .C1(n3238), .C2(n360), .A(n1061), 
        .ZN(n1059) );
  OAI221_X2 U365 ( .B1(n1062), .B2(n3274), .C1(n3309), .C2(n47), .A(n1063), 
        .ZN(n2642) );
  AOI221_X2 U368 ( .B1(ymem_data2[139]), .B2(n3277), .C1(ymem_data2[203]), 
        .C2(n3296), .A(n1069), .ZN(n1068) );
  OAI22_X2 U369 ( .A1(n3305), .A2(n551), .B1(n3303), .B2(n615), .ZN(n1069) );
  AOI221_X2 U370 ( .B1(ymem_data1[139]), .B2(n3292), .C1(ymem_data1[203]), 
        .C2(n3257), .A(n1070), .ZN(n1067) );
  OAI22_X2 U371 ( .A1(n3307), .A2(n359), .B1(n3284), .B2(n423), .ZN(n1070) );
  AOI221_X2 U373 ( .B1(ymem_data2[139]), .B2(n3271), .C1(ymem_data2[203]), 
        .C2(n3268), .A(n1073), .ZN(n1072) );
  OAI22_X2 U374 ( .A1(n3266), .A2(n551), .B1(n3264), .B2(n615), .ZN(n1073) );
  AOI221_X2 U375 ( .B1(ymem_data1[11]), .B2(n3263), .C1(ymem_data1[75]), .C2(
        n854), .A(n1074), .ZN(n1071) );
  OAI22_X2 U376 ( .A1(n856), .A2(n231), .B1(n3255), .B2(n295), .ZN(n1074) );
  AOI221_X2 U378 ( .B1(ymem_data1[11]), .B2(n3293), .C1(ymem_data2[203]), .C2(
        n860), .A(n1077), .ZN(n1076) );
  OAI22_X2 U379 ( .A1(n862), .A2(n359), .B1(n3249), .B2(n295), .ZN(n1077) );
  OAI22_X2 U382 ( .A1(n3240), .A2(n551), .B1(n99), .B2(n487), .ZN(n1079) );
  OAI221_X2 U383 ( .B1(n3249), .B2(n295), .C1(n3238), .C2(n359), .A(n1080), 
        .ZN(n1078) );
  OAI221_X2 U385 ( .B1(n1081), .B2(n3275), .C1(n3309), .C2(n46), .A(n1082), 
        .ZN(n2643) );
  AOI221_X2 U388 ( .B1(ymem_data2[140]), .B2(n3277), .C1(ymem_data2[204]), 
        .C2(n3296), .A(n1088), .ZN(n1087) );
  OAI22_X2 U389 ( .A1(n3305), .A2(n550), .B1(n3303), .B2(n614), .ZN(n1088) );
  AOI221_X2 U390 ( .B1(ymem_data1[140]), .B2(n110), .C1(ymem_data1[204]), .C2(
        n3258), .A(n1089), .ZN(n1086) );
  OAI22_X2 U394 ( .A1(n3266), .A2(n550), .B1(n3264), .B2(n614), .ZN(n1092) );
  AOI221_X2 U395 ( .B1(ymem_data1[12]), .B2(n3262), .C1(ymem_data1[76]), .C2(
        n854), .A(n1093), .ZN(n1090) );
  OAI22_X2 U396 ( .A1(n3259), .A2(n230), .B1(n3255), .B2(n294), .ZN(n1093) );
  AOI221_X2 U398 ( .B1(ymem_data1[12]), .B2(n3294), .C1(ymem_data2[204]), .C2(
        n860), .A(n1096), .ZN(n1095) );
  OAI22_X2 U399 ( .A1(n862), .A2(n358), .B1(n3249), .B2(n294), .ZN(n1096) );
  OAI22_X2 U402 ( .A1(n869), .A2(n550), .B1(n99), .B2(n486), .ZN(n1098) );
  OAI221_X2 U403 ( .B1(n863), .B2(n294), .C1(n3238), .C2(n358), .A(n1099), 
        .ZN(n1097) );
  OAI221_X2 U405 ( .B1(n1100), .B2(n3274), .C1(n3309), .C2(n45), .A(n1101), 
        .ZN(n2644) );
  AOI221_X2 U408 ( .B1(ymem_data2[141]), .B2(n3277), .C1(ymem_data2[205]), 
        .C2(n3296), .A(n1107), .ZN(n1106) );
  OAI22_X2 U409 ( .A1(n3305), .A2(n549), .B1(n3303), .B2(n613), .ZN(n1107) );
  AOI221_X2 U410 ( .B1(ymem_data1[141]), .B2(n110), .C1(ymem_data1[205]), .C2(
        n3257), .A(n1108), .ZN(n1105) );
  OAI22_X2 U411 ( .A1(n3307), .A2(n357), .B1(n778), .B2(n421), .ZN(n1108) );
  OAI22_X2 U414 ( .A1(n3266), .A2(n549), .B1(n3264), .B2(n613), .ZN(n1111) );
  AOI221_X2 U415 ( .B1(ymem_data1[13]), .B2(n3262), .C1(ymem_data1[77]), .C2(
        n854), .A(n1112), .ZN(n1109) );
  OAI22_X2 U416 ( .A1(n856), .A2(n229), .B1(n3255), .B2(n293), .ZN(n1112) );
  AOI221_X2 U418 ( .B1(ymem_data1[13]), .B2(n3294), .C1(ymem_data2[205]), .C2(
        n3253), .A(n1115), .ZN(n1114) );
  OAI22_X2 U422 ( .A1(n3240), .A2(n549), .B1(n99), .B2(n485), .ZN(n1117) );
  OAI221_X2 U425 ( .B1(n1119), .B2(n3275), .C1(n3309), .C2(n44), .A(n1120), 
        .ZN(n2645) );
  AOI221_X2 U428 ( .B1(ymem_data2[142]), .B2(n3277), .C1(ymem_data2[206]), 
        .C2(n3296), .A(n1126), .ZN(n1125) );
  OAI22_X2 U429 ( .A1(n3305), .A2(n548), .B1(n3303), .B2(n612), .ZN(n1126) );
  AOI221_X2 U430 ( .B1(ymem_data1[142]), .B2(n110), .C1(ymem_data1[206]), .C2(
        n3257), .A(n1127), .ZN(n1124) );
  OAI22_X2 U431 ( .A1(n3307), .A2(n356), .B1(n778), .B2(n420), .ZN(n1127) );
  AOI221_X2 U433 ( .B1(ymem_data2[142]), .B2(n3271), .C1(ymem_data2[206]), 
        .C2(n849), .A(n1130), .ZN(n1129) );
  OAI22_X2 U434 ( .A1(n3266), .A2(n548), .B1(n3264), .B2(n612), .ZN(n1130) );
  AOI221_X2 U435 ( .B1(ymem_data1[14]), .B2(n3262), .C1(ymem_data1[78]), .C2(
        n854), .A(n1131), .ZN(n1128) );
  OAI22_X2 U436 ( .A1(n856), .A2(n228), .B1(n3255), .B2(n292), .ZN(n1131) );
  AOI221_X2 U438 ( .B1(ymem_data1[14]), .B2(n3294), .C1(ymem_data2[206]), .C2(
        n3253), .A(n1134), .ZN(n1133) );
  OAI22_X2 U442 ( .A1(n3240), .A2(n548), .B1(n99), .B2(n484), .ZN(n1136) );
  OAI221_X2 U445 ( .B1(n1138), .B2(n3274), .C1(n3309), .C2(n43), .A(n1139), 
        .ZN(n2646) );
  AOI221_X2 U448 ( .B1(ymem_data2[143]), .B2(n3277), .C1(ymem_data2[207]), 
        .C2(n3296), .A(n1145), .ZN(n1144) );
  OAI22_X2 U449 ( .A1(n3305), .A2(n547), .B1(n3303), .B2(n611), .ZN(n1145) );
  AOI221_X2 U450 ( .B1(ymem_data1[143]), .B2(n110), .C1(ymem_data1[207]), .C2(
        n3257), .A(n1146), .ZN(n1143) );
  OAI22_X2 U451 ( .A1(n3307), .A2(n355), .B1(n778), .B2(n419), .ZN(n1146) );
  AOI221_X2 U453 ( .B1(ymem_data2[143]), .B2(n3271), .C1(ymem_data2[207]), 
        .C2(n849), .A(n1149), .ZN(n1148) );
  OAI22_X2 U454 ( .A1(n3266), .A2(n547), .B1(n3264), .B2(n611), .ZN(n1149) );
  AOI221_X2 U455 ( .B1(ymem_data1[15]), .B2(n3262), .C1(ymem_data1[79]), .C2(
        n854), .A(n1150), .ZN(n1147) );
  OAI22_X2 U456 ( .A1(n856), .A2(n227), .B1(n3255), .B2(n291), .ZN(n1150) );
  AOI221_X2 U458 ( .B1(ymem_data1[15]), .B2(n3294), .C1(ymem_data2[207]), .C2(
        n3253), .A(n1153), .ZN(n1152) );
  OAI22_X2 U462 ( .A1(n3240), .A2(n547), .B1(n99), .B2(n483), .ZN(n1155) );
  OAI221_X2 U463 ( .B1(n3249), .B2(n291), .C1(n870), .C2(n355), .A(n1156), 
        .ZN(n1154) );
  OAI221_X2 U465 ( .B1(n1157), .B2(n3275), .C1(n3309), .C2(n42), .A(n1158), 
        .ZN(n2647) );
  AOI221_X2 U468 ( .B1(ymem_data2[144]), .B2(n3277), .C1(ymem_data2[208]), 
        .C2(n3296), .A(n1164), .ZN(n1163) );
  OAI22_X2 U469 ( .A1(n3305), .A2(n546), .B1(n3303), .B2(n610), .ZN(n1164) );
  AOI221_X2 U470 ( .B1(ymem_data1[144]), .B2(n110), .C1(ymem_data1[208]), .C2(
        n3257), .A(n1165), .ZN(n1162) );
  OAI22_X2 U471 ( .A1(n3307), .A2(n354), .B1(n778), .B2(n418), .ZN(n1165) );
  AOI221_X2 U473 ( .B1(ymem_data2[144]), .B2(n3271), .C1(ymem_data2[208]), 
        .C2(n849), .A(n1168), .ZN(n1167) );
  OAI22_X2 U474 ( .A1(n3266), .A2(n546), .B1(n3264), .B2(n610), .ZN(n1168) );
  AOI221_X2 U475 ( .B1(ymem_data1[16]), .B2(n3262), .C1(ymem_data1[80]), .C2(
        n854), .A(n1169), .ZN(n1166) );
  OAI22_X2 U476 ( .A1(n856), .A2(n226), .B1(n3255), .B2(n290), .ZN(n1169) );
  AOI221_X2 U478 ( .B1(ymem_data1[16]), .B2(n3293), .C1(ymem_data2[208]), .C2(
        n3253), .A(n1172), .ZN(n1171) );
  OAI22_X2 U479 ( .A1(n862), .A2(n354), .B1(n3249), .B2(n290), .ZN(n1172) );
  OAI22_X2 U482 ( .A1(n3240), .A2(n546), .B1(n99), .B2(n482), .ZN(n1174) );
  OAI221_X2 U483 ( .B1(n3249), .B2(n290), .C1(n870), .C2(n354), .A(n1175), 
        .ZN(n1173) );
  OAI221_X2 U485 ( .B1(n1176), .B2(n3274), .C1(n3309), .C2(n41), .A(n1177), 
        .ZN(n2648) );
  AOI221_X2 U488 ( .B1(ymem_data2[145]), .B2(n3277), .C1(ymem_data2[209]), 
        .C2(n3296), .A(n1183), .ZN(n1182) );
  OAI22_X2 U489 ( .A1(n3305), .A2(n545), .B1(n3303), .B2(n609), .ZN(n1183) );
  AOI221_X2 U490 ( .B1(ymem_data1[145]), .B2(n110), .C1(ymem_data1[209]), .C2(
        n3257), .A(n1184), .ZN(n1181) );
  OAI22_X2 U491 ( .A1(n3307), .A2(n353), .B1(n778), .B2(n417), .ZN(n1184) );
  AOI221_X2 U493 ( .B1(ymem_data2[145]), .B2(n3271), .C1(ymem_data2[209]), 
        .C2(n849), .A(n1187), .ZN(n1186) );
  OAI22_X2 U494 ( .A1(n3266), .A2(n545), .B1(n3264), .B2(n609), .ZN(n1187) );
  AOI221_X2 U495 ( .B1(ymem_data1[17]), .B2(n3262), .C1(ymem_data1[81]), .C2(
        n854), .A(n1188), .ZN(n1185) );
  OAI22_X2 U496 ( .A1(n856), .A2(n225), .B1(n3255), .B2(n289), .ZN(n1188) );
  AOI221_X2 U498 ( .B1(ymem_data1[17]), .B2(n3294), .C1(ymem_data2[209]), .C2(
        n860), .A(n1191), .ZN(n1190) );
  OAI22_X2 U499 ( .A1(n862), .A2(n353), .B1(n3249), .B2(n289), .ZN(n1191) );
  OAI22_X2 U502 ( .A1(n869), .A2(n545), .B1(n99), .B2(n481), .ZN(n1193) );
  OAI221_X2 U503 ( .B1(n3249), .B2(n289), .C1(n870), .C2(n353), .A(n1194), 
        .ZN(n1192) );
  OAI221_X2 U505 ( .B1(n1195), .B2(n3275), .C1(n3309), .C2(n40), .A(n1196), 
        .ZN(n2649) );
  AOI221_X2 U508 ( .B1(ymem_data2[146]), .B2(n3277), .C1(ymem_data2[210]), 
        .C2(n3296), .A(n1202), .ZN(n1201) );
  OAI22_X2 U509 ( .A1(n3305), .A2(n544), .B1(n3303), .B2(n608), .ZN(n1202) );
  AOI221_X2 U510 ( .B1(ymem_data1[146]), .B2(n110), .C1(ymem_data1[210]), .C2(
        n3257), .A(n1203), .ZN(n1200) );
  OAI22_X2 U511 ( .A1(n3307), .A2(n352), .B1(n778), .B2(n416), .ZN(n1203) );
  AOI221_X2 U513 ( .B1(ymem_data2[146]), .B2(n3271), .C1(ymem_data2[210]), 
        .C2(n3268), .A(n1206), .ZN(n1205) );
  OAI22_X2 U514 ( .A1(n3266), .A2(n544), .B1(n3264), .B2(n608), .ZN(n1206) );
  AOI221_X2 U515 ( .B1(ymem_data1[18]), .B2(n3262), .C1(ymem_data1[82]), .C2(
        n854), .A(n1207), .ZN(n1204) );
  OAI22_X2 U516 ( .A1(n856), .A2(n224), .B1(n3255), .B2(n288), .ZN(n1207) );
  AOI221_X2 U518 ( .B1(ymem_data1[18]), .B2(n3293), .C1(ymem_data2[210]), .C2(
        n3253), .A(n1210), .ZN(n1209) );
  OAI22_X2 U519 ( .A1(n862), .A2(n352), .B1(n3249), .B2(n288), .ZN(n1210) );
  OAI22_X2 U522 ( .A1(n869), .A2(n544), .B1(n99), .B2(n480), .ZN(n1212) );
  OAI221_X2 U523 ( .B1(n863), .B2(n288), .C1(n870), .C2(n352), .A(n1213), .ZN(
        n1211) );
  OAI221_X2 U525 ( .B1(n1214), .B2(n3274), .C1(n3309), .C2(n39), .A(n1215), 
        .ZN(n2650) );
  AOI221_X2 U528 ( .B1(ymem_data2[147]), .B2(n3277), .C1(ymem_data2[211]), 
        .C2(n3296), .A(n1221), .ZN(n1220) );
  OAI22_X2 U529 ( .A1(n3305), .A2(n543), .B1(n3303), .B2(n607), .ZN(n1221) );
  AOI221_X2 U530 ( .B1(ymem_data1[147]), .B2(n110), .C1(ymem_data1[211]), .C2(
        n3257), .A(n1222), .ZN(n1219) );
  OAI22_X2 U531 ( .A1(n3307), .A2(n351), .B1(n778), .B2(n415), .ZN(n1222) );
  AOI221_X2 U533 ( .B1(ymem_data2[147]), .B2(n3271), .C1(ymem_data2[211]), 
        .C2(n3268), .A(n1225), .ZN(n1224) );
  OAI22_X2 U534 ( .A1(n3266), .A2(n543), .B1(n3264), .B2(n607), .ZN(n1225) );
  AOI221_X2 U535 ( .B1(ymem_data1[19]), .B2(n3262), .C1(ymem_data1[83]), .C2(
        n854), .A(n1226), .ZN(n1223) );
  OAI22_X2 U536 ( .A1(n856), .A2(n223), .B1(n3255), .B2(n287), .ZN(n1226) );
  AOI221_X2 U538 ( .B1(ymem_data1[19]), .B2(n3294), .C1(ymem_data2[211]), .C2(
        n860), .A(n1229), .ZN(n1228) );
  OAI22_X2 U539 ( .A1(n3251), .A2(n351), .B1(n3248), .B2(n287), .ZN(n1229) );
  OAI22_X2 U542 ( .A1(n869), .A2(n543), .B1(n99), .B2(n479), .ZN(n1231) );
  OAI221_X2 U543 ( .B1(n3249), .B2(n287), .C1(n870), .C2(n351), .A(n1232), 
        .ZN(n1230) );
  OAI221_X2 U545 ( .B1(n1233), .B2(n3275), .C1(n3309), .C2(n38), .A(n1234), 
        .ZN(n2651) );
  AOI221_X2 U548 ( .B1(ymem_data2[148]), .B2(n3277), .C1(ymem_data2[212]), 
        .C2(n3296), .A(n1240), .ZN(n1239) );
  OAI22_X2 U549 ( .A1(n3305), .A2(n542), .B1(n3303), .B2(n606), .ZN(n1240) );
  AOI221_X2 U550 ( .B1(ymem_data1[148]), .B2(n110), .C1(ymem_data1[212]), .C2(
        n3257), .A(n1241), .ZN(n1238) );
  OAI22_X2 U551 ( .A1(n3307), .A2(n350), .B1(n778), .B2(n414), .ZN(n1241) );
  AOI221_X2 U553 ( .B1(ymem_data2[148]), .B2(n3271), .C1(ymem_data2[212]), 
        .C2(n3268), .A(n1244), .ZN(n1243) );
  OAI22_X2 U554 ( .A1(n3266), .A2(n542), .B1(n3264), .B2(n606), .ZN(n1244) );
  AOI221_X2 U555 ( .B1(ymem_data1[20]), .B2(n3262), .C1(ymem_data1[84]), .C2(
        n854), .A(n1245), .ZN(n1242) );
  OAI22_X2 U556 ( .A1(n856), .A2(n222), .B1(n3255), .B2(n286), .ZN(n1245) );
  AOI221_X2 U558 ( .B1(ymem_data1[20]), .B2(n3293), .C1(ymem_data2[212]), .C2(
        n860), .A(n1248), .ZN(n1247) );
  OAI22_X2 U559 ( .A1(n3251), .A2(n350), .B1(n3248), .B2(n286), .ZN(n1248) );
  OAI22_X2 U562 ( .A1(n869), .A2(n542), .B1(n99), .B2(n478), .ZN(n1250) );
  OAI221_X2 U563 ( .B1(n3249), .B2(n286), .C1(n870), .C2(n350), .A(n1251), 
        .ZN(n1249) );
  OAI221_X2 U565 ( .B1(n1252), .B2(n3274), .C1(n3309), .C2(n37), .A(n1253), 
        .ZN(n2652) );
  AOI221_X2 U568 ( .B1(ymem_data2[149]), .B2(n3277), .C1(ymem_data2[213]), 
        .C2(n3296), .A(n1259), .ZN(n1258) );
  OAI22_X2 U569 ( .A1(n3305), .A2(n541), .B1(n3303), .B2(n605), .ZN(n1259) );
  AOI221_X2 U570 ( .B1(ymem_data1[149]), .B2(n110), .C1(ymem_data1[213]), .C2(
        n3257), .A(n1260), .ZN(n1257) );
  OAI22_X2 U571 ( .A1(n3307), .A2(n349), .B1(n778), .B2(n413), .ZN(n1260) );
  AOI221_X2 U573 ( .B1(ymem_data2[149]), .B2(n3271), .C1(ymem_data2[213]), 
        .C2(n3268), .A(n1263), .ZN(n1262) );
  OAI22_X2 U574 ( .A1(n3266), .A2(n541), .B1(n3264), .B2(n605), .ZN(n1263) );
  AOI221_X2 U575 ( .B1(ymem_data1[21]), .B2(n3262), .C1(ymem_data1[85]), .C2(
        n854), .A(n1264), .ZN(n1261) );
  OAI22_X2 U576 ( .A1(n856), .A2(n221), .B1(n3255), .B2(n285), .ZN(n1264) );
  AOI221_X2 U578 ( .B1(ymem_data1[21]), .B2(n3294), .C1(ymem_data2[213]), .C2(
        n860), .A(n1267), .ZN(n1266) );
  OAI22_X2 U579 ( .A1(n3251), .A2(n349), .B1(n3248), .B2(n285), .ZN(n1267) );
  OAI22_X2 U582 ( .A1(n869), .A2(n541), .B1(n99), .B2(n477), .ZN(n1269) );
  OAI221_X2 U583 ( .B1(n3249), .B2(n285), .C1(n870), .C2(n349), .A(n1270), 
        .ZN(n1268) );
  OAI221_X2 U585 ( .B1(n1271), .B2(n3275), .C1(n3309), .C2(n36), .A(n1272), 
        .ZN(n2653) );
  AOI221_X2 U588 ( .B1(ymem_data2[150]), .B2(n3276), .C1(ymem_data2[214]), 
        .C2(n3296), .A(n1278), .ZN(n1277) );
  OAI22_X2 U589 ( .A1(n3305), .A2(n540), .B1(n3303), .B2(n604), .ZN(n1278) );
  AOI221_X2 U590 ( .B1(ymem_data1[150]), .B2(n110), .C1(ymem_data1[214]), .C2(
        n3257), .A(n1279), .ZN(n1276) );
  OAI22_X2 U591 ( .A1(n3307), .A2(n348), .B1(n778), .B2(n412), .ZN(n1279) );
  AOI221_X2 U593 ( .B1(ymem_data2[150]), .B2(n3270), .C1(ymem_data2[214]), 
        .C2(n3268), .A(n1282), .ZN(n1281) );
  OAI22_X2 U594 ( .A1(n3266), .A2(n540), .B1(n3264), .B2(n604), .ZN(n1282) );
  AOI221_X2 U595 ( .B1(ymem_data1[22]), .B2(n3262), .C1(ymem_data1[86]), .C2(
        n3261), .A(n1283), .ZN(n1280) );
  AOI221_X2 U598 ( .B1(ymem_data1[22]), .B2(n3294), .C1(ymem_data2[214]), .C2(
        n3253), .A(n1286), .ZN(n1285) );
  OAI22_X2 U599 ( .A1(n3251), .A2(n348), .B1(n3248), .B2(n284), .ZN(n1286) );
  OAI22_X2 U602 ( .A1(n869), .A2(n540), .B1(n99), .B2(n476), .ZN(n1288) );
  OAI221_X2 U603 ( .B1(n3249), .B2(n284), .C1(n870), .C2(n348), .A(n1289), 
        .ZN(n1287) );
  OAI221_X2 U605 ( .B1(n1290), .B2(n3275), .C1(n3309), .C2(n35), .A(n1291), 
        .ZN(n2654) );
  AOI221_X2 U608 ( .B1(ymem_data2[151]), .B2(n3276), .C1(ymem_data2[215]), 
        .C2(n3297), .A(n1297), .ZN(n1296) );
  OAI22_X2 U609 ( .A1(n3305), .A2(n539), .B1(n3303), .B2(n603), .ZN(n1297) );
  AOI221_X2 U610 ( .B1(ymem_data1[151]), .B2(n110), .C1(ymem_data1[215]), .C2(
        n3257), .A(n1298), .ZN(n1295) );
  OAI22_X2 U611 ( .A1(n3307), .A2(n347), .B1(n778), .B2(n411), .ZN(n1298) );
  AOI221_X2 U613 ( .B1(ymem_data2[151]), .B2(n3270), .C1(ymem_data2[215]), 
        .C2(n3268), .A(n1301), .ZN(n1300) );
  OAI22_X2 U614 ( .A1(n3266), .A2(n539), .B1(n3264), .B2(n603), .ZN(n1301) );
  AOI221_X2 U615 ( .B1(ymem_data1[23]), .B2(n3262), .C1(ymem_data1[87]), .C2(
        n3261), .A(n1302), .ZN(n1299) );
  AOI221_X2 U618 ( .B1(ymem_data1[23]), .B2(n3294), .C1(ymem_data2[215]), .C2(
        n3253), .A(n1305), .ZN(n1304) );
  OAI22_X2 U619 ( .A1(n3251), .A2(n347), .B1(n3248), .B2(n283), .ZN(n1305) );
  OAI22_X2 U622 ( .A1(n869), .A2(n539), .B1(n99), .B2(n475), .ZN(n1307) );
  OAI221_X2 U623 ( .B1(n3248), .B2(n283), .C1(n3238), .C2(n347), .A(n1308), 
        .ZN(n1306) );
  OAI221_X2 U625 ( .B1(n1309), .B2(n3275), .C1(n3309), .C2(n34), .A(n1310), 
        .ZN(n2655) );
  AOI221_X2 U628 ( .B1(ymem_data2[152]), .B2(n3276), .C1(ymem_data2[216]), 
        .C2(n3296), .A(n1316), .ZN(n1315) );
  OAI22_X2 U629 ( .A1(n3305), .A2(n538), .B1(n3303), .B2(n602), .ZN(n1316) );
  AOI221_X2 U630 ( .B1(ymem_data1[152]), .B2(n3292), .C1(ymem_data1[216]), 
        .C2(n3257), .A(n1317), .ZN(n1314) );
  OAI22_X2 U631 ( .A1(n3307), .A2(n346), .B1(n3284), .B2(n410), .ZN(n1317) );
  AOI221_X2 U633 ( .B1(ymem_data2[152]), .B2(n3270), .C1(ymem_data2[216]), 
        .C2(n3268), .A(n1320), .ZN(n1319) );
  OAI22_X2 U634 ( .A1(n3266), .A2(n538), .B1(n3264), .B2(n602), .ZN(n1320) );
  AOI221_X2 U635 ( .B1(ymem_data1[24]), .B2(n3262), .C1(ymem_data1[88]), .C2(
        n3261), .A(n1321), .ZN(n1318) );
  AOI221_X2 U638 ( .B1(ymem_data1[24]), .B2(n3294), .C1(ymem_data2[216]), .C2(
        n860), .A(n1324), .ZN(n1323) );
  OAI22_X2 U642 ( .A1(n869), .A2(n538), .B1(n99), .B2(n474), .ZN(n1326) );
  OAI221_X2 U643 ( .B1(n3249), .B2(n282), .C1(n870), .C2(n346), .A(n1327), 
        .ZN(n1325) );
  OAI221_X2 U645 ( .B1(n1328), .B2(n3275), .C1(n3309), .C2(n33), .A(n1329), 
        .ZN(n2656) );
  AOI221_X2 U648 ( .B1(ymem_data2[153]), .B2(n3276), .C1(ymem_data2[217]), 
        .C2(n3297), .A(n1335), .ZN(n1334) );
  OAI22_X2 U649 ( .A1(n3305), .A2(n537), .B1(n3303), .B2(n601), .ZN(n1335) );
  AOI221_X2 U650 ( .B1(ymem_data1[153]), .B2(n3292), .C1(ymem_data1[217]), 
        .C2(n3257), .A(n1336), .ZN(n1333) );
  OAI22_X2 U651 ( .A1(n3307), .A2(n345), .B1(n3284), .B2(n409), .ZN(n1336) );
  AOI221_X2 U653 ( .B1(ymem_data2[153]), .B2(n3270), .C1(ymem_data2[217]), 
        .C2(n3268), .A(n1339), .ZN(n1338) );
  OAI22_X2 U654 ( .A1(n3266), .A2(n537), .B1(n3264), .B2(n601), .ZN(n1339) );
  AOI221_X2 U655 ( .B1(ymem_data1[25]), .B2(n3262), .C1(ymem_data1[89]), .C2(
        n3261), .A(n1340), .ZN(n1337) );
  AOI221_X2 U658 ( .B1(ymem_data1[25]), .B2(n3294), .C1(ymem_data2[217]), .C2(
        n860), .A(n1343), .ZN(n1342) );
  OAI22_X2 U662 ( .A1(n869), .A2(n537), .B1(n99), .B2(n473), .ZN(n1345) );
  OAI221_X2 U663 ( .B1(n3249), .B2(n281), .C1(n870), .C2(n345), .A(n1346), 
        .ZN(n1344) );
  OAI221_X2 U665 ( .B1(n1347), .B2(n3275), .C1(n3309), .C2(n32), .A(n1348), 
        .ZN(n2657) );
  AOI221_X2 U668 ( .B1(ymem_data2[154]), .B2(n3276), .C1(ymem_data2[218]), 
        .C2(n3296), .A(n1354), .ZN(n1353) );
  OAI22_X2 U669 ( .A1(n3305), .A2(n536), .B1(n3303), .B2(n600), .ZN(n1354) );
  AOI221_X2 U670 ( .B1(ymem_data1[154]), .B2(n110), .C1(ymem_data1[218]), .C2(
        n3257), .A(n1355), .ZN(n1352) );
  OAI22_X2 U671 ( .A1(n3307), .A2(n344), .B1(n3284), .B2(n408), .ZN(n1355) );
  AOI221_X2 U673 ( .B1(ymem_data2[154]), .B2(n3270), .C1(ymem_data2[218]), 
        .C2(n849), .A(n1358), .ZN(n1357) );
  OAI22_X2 U674 ( .A1(n3266), .A2(n536), .B1(n3264), .B2(n600), .ZN(n1358) );
  AOI221_X2 U675 ( .B1(ymem_data1[26]), .B2(n3263), .C1(ymem_data1[90]), .C2(
        n3261), .A(n1359), .ZN(n1356) );
  OAI22_X2 U676 ( .A1(n856), .A2(n216), .B1(n3255), .B2(n280), .ZN(n1359) );
  AOI221_X2 U678 ( .B1(ymem_data1[26]), .B2(n3294), .C1(ymem_data2[218]), .C2(
        n860), .A(n1362), .ZN(n1361) );
  OAI22_X2 U682 ( .A1(n869), .A2(n536), .B1(n99), .B2(n472), .ZN(n1364) );
  OAI221_X2 U683 ( .B1(n3249), .B2(n280), .C1(n3238), .C2(n344), .A(n1365), 
        .ZN(n1363) );
  OAI221_X2 U685 ( .B1(n1366), .B2(n3275), .C1(n3309), .C2(n31), .A(n1367), 
        .ZN(n2658) );
  AOI221_X2 U688 ( .B1(ymem_data2[155]), .B2(n3276), .C1(ymem_data2[219]), 
        .C2(n3297), .A(n1373), .ZN(n1372) );
  OAI22_X2 U689 ( .A1(n3305), .A2(n535), .B1(n3303), .B2(n599), .ZN(n1373) );
  AOI221_X2 U690 ( .B1(ymem_data1[155]), .B2(n3292), .C1(ymem_data1[219]), 
        .C2(n3257), .A(n1374), .ZN(n1371) );
  OAI22_X2 U691 ( .A1(n3307), .A2(n343), .B1(n3284), .B2(n407), .ZN(n1374) );
  AOI221_X2 U693 ( .B1(ymem_data2[155]), .B2(n3270), .C1(ymem_data2[219]), 
        .C2(n849), .A(n1377), .ZN(n1376) );
  OAI22_X2 U694 ( .A1(n3266), .A2(n535), .B1(n3264), .B2(n599), .ZN(n1377) );
  AOI221_X2 U695 ( .B1(ymem_data1[27]), .B2(n3263), .C1(ymem_data1[91]), .C2(
        n3261), .A(n1378), .ZN(n1375) );
  OAI22_X2 U696 ( .A1(n856), .A2(n215), .B1(n3255), .B2(n279), .ZN(n1378) );
  AOI221_X2 U698 ( .B1(ymem_data1[27]), .B2(n3294), .C1(ymem_data2[219]), .C2(
        n860), .A(n1381), .ZN(n1380) );
  OAI22_X2 U699 ( .A1(n862), .A2(n343), .B1(n863), .B2(n279), .ZN(n1381) );
  OAI22_X2 U702 ( .A1(n869), .A2(n535), .B1(n99), .B2(n471), .ZN(n1383) );
  OAI221_X2 U703 ( .B1(n863), .B2(n279), .C1(n3238), .C2(n343), .A(n1384), 
        .ZN(n1382) );
  OAI221_X2 U705 ( .B1(n1385), .B2(n3275), .C1(n3309), .C2(n30), .A(n1386), 
        .ZN(n2659) );
  AOI221_X2 U708 ( .B1(ymem_data2[156]), .B2(n3276), .C1(ymem_data2[220]), 
        .C2(n3296), .A(n1392), .ZN(n1391) );
  OAI22_X2 U709 ( .A1(n3305), .A2(n534), .B1(n3303), .B2(n598), .ZN(n1392) );
  AOI221_X2 U710 ( .B1(ymem_data1[156]), .B2(n110), .C1(ymem_data1[220]), .C2(
        n3258), .A(n1393), .ZN(n1390) );
  OAI22_X2 U711 ( .A1(n3307), .A2(n342), .B1(n3284), .B2(n406), .ZN(n1393) );
  AOI221_X2 U713 ( .B1(ymem_data2[156]), .B2(n3270), .C1(ymem_data2[220]), 
        .C2(n849), .A(n1396), .ZN(n1395) );
  OAI22_X2 U714 ( .A1(n3266), .A2(n534), .B1(n3264), .B2(n598), .ZN(n1396) );
  AOI221_X2 U715 ( .B1(ymem_data1[28]), .B2(n3263), .C1(ymem_data1[92]), .C2(
        n3261), .A(n1397), .ZN(n1394) );
  OAI22_X2 U716 ( .A1(n856), .A2(n214), .B1(n3255), .B2(n278), .ZN(n1397) );
  AOI221_X2 U718 ( .B1(ymem_data1[28]), .B2(n3294), .C1(ymem_data2[220]), .C2(
        n860), .A(n1400), .ZN(n1399) );
  OAI22_X2 U719 ( .A1(n862), .A2(n342), .B1(n3249), .B2(n278), .ZN(n1400) );
  OAI22_X2 U722 ( .A1(n869), .A2(n534), .B1(n99), .B2(n470), .ZN(n1402) );
  OAI221_X2 U723 ( .B1(n863), .B2(n278), .C1(n3238), .C2(n342), .A(n1403), 
        .ZN(n1401) );
  OAI221_X2 U725 ( .B1(n1404), .B2(n3275), .C1(n3309), .C2(n29), .A(n1405), 
        .ZN(n2660) );
  AOI221_X2 U728 ( .B1(ymem_data2[157]), .B2(n3276), .C1(ymem_data2[221]), 
        .C2(n3297), .A(n1411), .ZN(n1410) );
  OAI22_X2 U729 ( .A1(n3305), .A2(n533), .B1(n3303), .B2(n597), .ZN(n1411) );
  AOI221_X2 U730 ( .B1(ymem_data1[157]), .B2(n110), .C1(ymem_data1[221]), .C2(
        n3257), .A(n1412), .ZN(n1409) );
  OAI22_X2 U731 ( .A1(n3307), .A2(n341), .B1(n3284), .B2(n405), .ZN(n1412) );
  AOI221_X2 U733 ( .B1(ymem_data2[157]), .B2(n3270), .C1(ymem_data2[221]), 
        .C2(n849), .A(n1415), .ZN(n1414) );
  OAI22_X2 U734 ( .A1(n3266), .A2(n533), .B1(n3264), .B2(n597), .ZN(n1415) );
  AOI221_X2 U735 ( .B1(ymem_data1[29]), .B2(n3263), .C1(ymem_data1[93]), .C2(
        n854), .A(n1416), .ZN(n1413) );
  OAI22_X2 U736 ( .A1(n3259), .A2(n213), .B1(n857), .B2(n277), .ZN(n1416) );
  AOI221_X2 U738 ( .B1(ymem_data1[29]), .B2(n3294), .C1(ymem_data2[221]), .C2(
        n3253), .A(n1419), .ZN(n1418) );
  OAI22_X2 U742 ( .A1(n3240), .A2(n533), .B1(n99), .B2(n469), .ZN(n1421) );
  OAI221_X2 U743 ( .B1(n863), .B2(n277), .C1(n3238), .C2(n341), .A(n1422), 
        .ZN(n1420) );
  OAI221_X2 U745 ( .B1(n1423), .B2(n3275), .C1(n3309), .C2(n28), .A(n1424), 
        .ZN(n2661) );
  AOI221_X2 U748 ( .B1(ymem_data2[158]), .B2(n3276), .C1(ymem_data2[222]), 
        .C2(n3296), .A(n1430), .ZN(n1429) );
  OAI22_X2 U749 ( .A1(n3305), .A2(n532), .B1(n3303), .B2(n596), .ZN(n1430) );
  AOI221_X2 U750 ( .B1(ymem_data1[158]), .B2(n3292), .C1(ymem_data1[222]), 
        .C2(n3257), .A(n1431), .ZN(n1428) );
  OAI22_X2 U751 ( .A1(n3307), .A2(n340), .B1(n3284), .B2(n404), .ZN(n1431) );
  AOI221_X2 U753 ( .B1(ymem_data2[158]), .B2(n3270), .C1(ymem_data2[222]), 
        .C2(n849), .A(n1434), .ZN(n1433) );
  OAI22_X2 U754 ( .A1(n3266), .A2(n532), .B1(n3264), .B2(n596), .ZN(n1434) );
  AOI221_X2 U755 ( .B1(ymem_data1[30]), .B2(n3263), .C1(ymem_data1[94]), .C2(
        n854), .A(n1435), .ZN(n1432) );
  OAI22_X2 U756 ( .A1(n3259), .A2(n212), .B1(n857), .B2(n276), .ZN(n1435) );
  AOI221_X2 U758 ( .B1(ymem_data1[30]), .B2(n3294), .C1(ymem_data2[222]), .C2(
        n3253), .A(n1438), .ZN(n1437) );
  OAI22_X2 U762 ( .A1(n3240), .A2(n532), .B1(n99), .B2(n468), .ZN(n1440) );
  OAI221_X2 U763 ( .B1(n863), .B2(n276), .C1(n3238), .C2(n340), .A(n1441), 
        .ZN(n1439) );
  OAI221_X2 U765 ( .B1(n1442), .B2(n3275), .C1(n3309), .C2(n27), .A(n1443), 
        .ZN(n2662) );
  AOI221_X2 U768 ( .B1(ymem_data2[159]), .B2(n3276), .C1(ymem_data2[223]), 
        .C2(n3297), .A(n1449), .ZN(n1448) );
  OAI22_X2 U769 ( .A1(n3305), .A2(n531), .B1(n3303), .B2(n595), .ZN(n1449) );
  AOI221_X2 U770 ( .B1(ymem_data1[159]), .B2(n110), .C1(ymem_data1[223]), .C2(
        n3257), .A(n1450), .ZN(n1447) );
  OAI22_X2 U771 ( .A1(n3307), .A2(n339), .B1(n3284), .B2(n403), .ZN(n1450) );
  AOI221_X2 U773 ( .B1(ymem_data2[159]), .B2(n3270), .C1(ymem_data2[223]), 
        .C2(n849), .A(n1453), .ZN(n1452) );
  OAI22_X2 U774 ( .A1(n3266), .A2(n531), .B1(n3264), .B2(n595), .ZN(n1453) );
  AOI221_X2 U775 ( .B1(ymem_data1[31]), .B2(n3263), .C1(ymem_data1[95]), .C2(
        n854), .A(n1454), .ZN(n1451) );
  OAI22_X2 U776 ( .A1(n3259), .A2(n211), .B1(n3255), .B2(n275), .ZN(n1454) );
  AOI221_X2 U778 ( .B1(ymem_data1[31]), .B2(n3294), .C1(ymem_data2[223]), .C2(
        n3253), .A(n1457), .ZN(n1456) );
  OAI22_X2 U782 ( .A1(n3240), .A2(n531), .B1(n99), .B2(n467), .ZN(n1459) );
  OAI221_X2 U783 ( .B1(n3248), .B2(n275), .C1(n3238), .C2(n339), .A(n1460), 
        .ZN(n1458) );
  OAI221_X2 U785 ( .B1(n1461), .B2(n3275), .C1(n3309), .C2(n26), .A(n1462), 
        .ZN(n2663) );
  AOI221_X2 U788 ( .B1(ymem_data2[160]), .B2(n3276), .C1(ymem_data2[224]), 
        .C2(n3296), .A(n1468), .ZN(n1467) );
  OAI22_X2 U789 ( .A1(n3305), .A2(n530), .B1(n3303), .B2(n594), .ZN(n1468) );
  AOI221_X2 U790 ( .B1(ymem_data1[160]), .B2(n3292), .C1(ymem_data1[224]), 
        .C2(n3257), .A(n1469), .ZN(n1466) );
  OAI22_X2 U791 ( .A1(n3307), .A2(n338), .B1(n3284), .B2(n402), .ZN(n1469) );
  AOI221_X2 U793 ( .B1(ymem_data2[160]), .B2(n3270), .C1(ymem_data2[224]), 
        .C2(n849), .A(n1472), .ZN(n1471) );
  OAI22_X2 U794 ( .A1(n3266), .A2(n530), .B1(n3264), .B2(n594), .ZN(n1472) );
  AOI221_X2 U795 ( .B1(ymem_data1[32]), .B2(n3263), .C1(ymem_data1[96]), .C2(
        n854), .A(n1473), .ZN(n1470) );
  OAI22_X2 U796 ( .A1(n3259), .A2(n210), .B1(n3255), .B2(n274), .ZN(n1473) );
  AOI221_X2 U798 ( .B1(ymem_data1[32]), .B2(n3294), .C1(ymem_data2[224]), .C2(
        n3253), .A(n1476), .ZN(n1475) );
  OAI22_X2 U799 ( .A1(n862), .A2(n338), .B1(n3249), .B2(n274), .ZN(n1476) );
  OAI22_X2 U802 ( .A1(n3240), .A2(n530), .B1(n99), .B2(n466), .ZN(n1478) );
  OAI221_X2 U803 ( .B1(n863), .B2(n274), .C1(n3238), .C2(n338), .A(n1479), 
        .ZN(n1477) );
  OAI221_X2 U805 ( .B1(n1480), .B2(n3275), .C1(n3309), .C2(n25), .A(n1481), 
        .ZN(n2664) );
  AOI221_X2 U808 ( .B1(ymem_data2[161]), .B2(n3276), .C1(ymem_data2[225]), 
        .C2(n3297), .A(n1487), .ZN(n1486) );
  OAI22_X2 U809 ( .A1(n3305), .A2(n529), .B1(n3303), .B2(n593), .ZN(n1487) );
  AOI221_X2 U810 ( .B1(ymem_data1[161]), .B2(n110), .C1(ymem_data1[225]), .C2(
        n3257), .A(n1488), .ZN(n1485) );
  OAI22_X2 U811 ( .A1(n3307), .A2(n337), .B1(n3284), .B2(n401), .ZN(n1488) );
  AOI221_X2 U813 ( .B1(ymem_data2[161]), .B2(n3270), .C1(ymem_data2[225]), 
        .C2(n849), .A(n1491), .ZN(n1490) );
  OAI22_X2 U814 ( .A1(n3266), .A2(n529), .B1(n3264), .B2(n593), .ZN(n1491) );
  AOI221_X2 U815 ( .B1(ymem_data1[33]), .B2(n3263), .C1(ymem_data1[97]), .C2(
        n3261), .A(n1492), .ZN(n1489) );
  OAI22_X2 U816 ( .A1(n3259), .A2(n209), .B1(n3255), .B2(n273), .ZN(n1492) );
  AOI221_X2 U818 ( .B1(ymem_data1[33]), .B2(n3294), .C1(ymem_data2[225]), .C2(
        n3253), .A(n1495), .ZN(n1494) );
  OAI22_X2 U819 ( .A1(n862), .A2(n337), .B1(n3248), .B2(n273), .ZN(n1495) );
  OAI22_X2 U822 ( .A1(n3240), .A2(n529), .B1(n99), .B2(n465), .ZN(n1497) );
  OAI221_X2 U823 ( .B1(n863), .B2(n273), .C1(n3238), .C2(n337), .A(n1498), 
        .ZN(n1496) );
  OAI221_X2 U825 ( .B1(n1499), .B2(n3275), .C1(n3309), .C2(n24), .A(n1500), 
        .ZN(n2665) );
  AOI221_X2 U828 ( .B1(ymem_data2[162]), .B2(n3276), .C1(ymem_data2[226]), 
        .C2(n3296), .A(n1506), .ZN(n1505) );
  OAI22_X2 U829 ( .A1(n3305), .A2(n528), .B1(n3303), .B2(n592), .ZN(n1506) );
  AOI221_X2 U830 ( .B1(ymem_data1[162]), .B2(n3292), .C1(ymem_data1[226]), 
        .C2(n3257), .A(n1507), .ZN(n1504) );
  OAI22_X2 U831 ( .A1(n3307), .A2(n336), .B1(n3284), .B2(n400), .ZN(n1507) );
  AOI221_X2 U833 ( .B1(ymem_data2[162]), .B2(n3270), .C1(ymem_data2[226]), 
        .C2(n849), .A(n1510), .ZN(n1509) );
  OAI22_X2 U834 ( .A1(n3266), .A2(n528), .B1(n3264), .B2(n592), .ZN(n1510) );
  AOI221_X2 U835 ( .B1(ymem_data1[34]), .B2(n3263), .C1(ymem_data1[98]), .C2(
        n3261), .A(n1511), .ZN(n1508) );
  OAI22_X2 U836 ( .A1(n3259), .A2(n208), .B1(n3255), .B2(n272), .ZN(n1511) );
  AOI221_X2 U838 ( .B1(ymem_data1[34]), .B2(n3294), .C1(ymem_data2[226]), .C2(
        n3253), .A(n1514), .ZN(n1513) );
  OAI22_X2 U842 ( .A1(n3240), .A2(n528), .B1(n99), .B2(n464), .ZN(n1516) );
  OAI221_X2 U843 ( .B1(n3248), .B2(n272), .C1(n3238), .C2(n336), .A(n1517), 
        .ZN(n1515) );
  OAI221_X2 U845 ( .B1(n1518), .B2(n3274), .C1(n3309), .C2(n23), .A(n1519), 
        .ZN(n2666) );
  AOI221_X2 U848 ( .B1(ymem_data2[163]), .B2(n3276), .C1(ymem_data2[227]), 
        .C2(n3297), .A(n1525), .ZN(n1524) );
  OAI22_X2 U849 ( .A1(n3305), .A2(n527), .B1(n3303), .B2(n591), .ZN(n1525) );
  AOI221_X2 U850 ( .B1(ymem_data1[163]), .B2(n3292), .C1(ymem_data1[227]), 
        .C2(n3257), .A(n1526), .ZN(n1523) );
  OAI22_X2 U851 ( .A1(n3307), .A2(n335), .B1(n3284), .B2(n399), .ZN(n1526) );
  AOI221_X2 U853 ( .B1(ymem_data2[163]), .B2(n3270), .C1(ymem_data2[227]), 
        .C2(n849), .A(n1529), .ZN(n1528) );
  OAI22_X2 U854 ( .A1(n3266), .A2(n527), .B1(n3264), .B2(n591), .ZN(n1529) );
  AOI221_X2 U855 ( .B1(ymem_data1[35]), .B2(n3263), .C1(ymem_data1[99]), .C2(
        n3261), .A(n1530), .ZN(n1527) );
  OAI22_X2 U856 ( .A1(n3259), .A2(n207), .B1(n3255), .B2(n271), .ZN(n1530) );
  AOI221_X2 U858 ( .B1(ymem_data1[35]), .B2(n3293), .C1(ymem_data2[227]), .C2(
        n3253), .A(n1533), .ZN(n1532) );
  OAI22_X2 U859 ( .A1(n862), .A2(n335), .B1(n3248), .B2(n271), .ZN(n1533) );
  OAI22_X2 U862 ( .A1(n3240), .A2(n527), .B1(n99), .B2(n463), .ZN(n1535) );
  OAI221_X2 U863 ( .B1(n863), .B2(n271), .C1(n3238), .C2(n335), .A(n1536), 
        .ZN(n1534) );
  OAI221_X2 U865 ( .B1(n1537), .B2(n3274), .C1(n3309), .C2(n22), .A(n1538), 
        .ZN(n2667) );
  AOI221_X2 U868 ( .B1(ymem_data2[164]), .B2(n3277), .C1(ymem_data2[228]), 
        .C2(n3297), .A(n1544), .ZN(n1543) );
  OAI22_X2 U869 ( .A1(n3305), .A2(n526), .B1(n3303), .B2(n590), .ZN(n1544) );
  AOI221_X2 U870 ( .B1(ymem_data1[164]), .B2(n3292), .C1(ymem_data1[228]), 
        .C2(n3257), .A(n1545), .ZN(n1542) );
  OAI22_X2 U871 ( .A1(n3307), .A2(n334), .B1(n3284), .B2(n398), .ZN(n1545) );
  AOI221_X2 U873 ( .B1(ymem_data2[164]), .B2(n3271), .C1(ymem_data2[228]), 
        .C2(n849), .A(n1548), .ZN(n1547) );
  OAI22_X2 U874 ( .A1(n3266), .A2(n526), .B1(n3264), .B2(n590), .ZN(n1548) );
  AOI221_X2 U875 ( .B1(ymem_data1[36]), .B2(n3263), .C1(ymem_data1[100]), .C2(
        n854), .A(n1549), .ZN(n1546) );
  OAI22_X2 U876 ( .A1(n3259), .A2(n206), .B1(n3255), .B2(n270), .ZN(n1549) );
  AOI221_X2 U878 ( .B1(ymem_data1[36]), .B2(n3293), .C1(ymem_data2[228]), .C2(
        n3253), .A(n1552), .ZN(n1551) );
  OAI22_X2 U879 ( .A1(n3251), .A2(n334), .B1(n3249), .B2(n270), .ZN(n1552) );
  OAI22_X2 U882 ( .A1(n3240), .A2(n526), .B1(n99), .B2(n462), .ZN(n1554) );
  OAI221_X2 U883 ( .B1(n3249), .B2(n270), .C1(n3238), .C2(n334), .A(n1555), 
        .ZN(n1553) );
  OAI221_X2 U885 ( .B1(n1556), .B2(n3274), .C1(n3309), .C2(n21), .A(n1557), 
        .ZN(n2668) );
  AOI221_X2 U888 ( .B1(ymem_data2[165]), .B2(n3276), .C1(ymem_data2[229]), 
        .C2(n3297), .A(n1563), .ZN(n1562) );
  OAI22_X2 U889 ( .A1(n3305), .A2(n525), .B1(n3303), .B2(n589), .ZN(n1563) );
  AOI221_X2 U890 ( .B1(ymem_data1[165]), .B2(n3292), .C1(ymem_data1[229]), 
        .C2(n3257), .A(n1564), .ZN(n1561) );
  OAI22_X2 U891 ( .A1(n3307), .A2(n333), .B1(n3284), .B2(n397), .ZN(n1564) );
  AOI221_X2 U893 ( .B1(ymem_data2[165]), .B2(n3270), .C1(ymem_data2[229]), 
        .C2(n849), .A(n1567), .ZN(n1566) );
  OAI22_X2 U894 ( .A1(n3266), .A2(n525), .B1(n3264), .B2(n589), .ZN(n1567) );
  AOI221_X2 U895 ( .B1(ymem_data1[37]), .B2(n3263), .C1(ymem_data1[101]), .C2(
        n3261), .A(n1568), .ZN(n1565) );
  OAI22_X2 U896 ( .A1(n3259), .A2(n205), .B1(n3255), .B2(n269), .ZN(n1568) );
  AOI221_X2 U898 ( .B1(ymem_data1[37]), .B2(n3293), .C1(ymem_data2[229]), .C2(
        n3253), .A(n1571), .ZN(n1570) );
  OAI22_X2 U899 ( .A1(n3251), .A2(n333), .B1(n3248), .B2(n269), .ZN(n1571) );
  OAI22_X2 U902 ( .A1(n3240), .A2(n525), .B1(n99), .B2(n461), .ZN(n1573) );
  OAI221_X2 U903 ( .B1(n3248), .B2(n269), .C1(n3238), .C2(n333), .A(n1574), 
        .ZN(n1572) );
  OAI221_X2 U905 ( .B1(n1575), .B2(n3274), .C1(n3309), .C2(n20), .A(n1576), 
        .ZN(n2669) );
  AOI221_X2 U908 ( .B1(ymem_data2[166]), .B2(n3277), .C1(ymem_data2[230]), 
        .C2(n3297), .A(n1582), .ZN(n1581) );
  OAI22_X2 U909 ( .A1(n3305), .A2(n524), .B1(n3303), .B2(n588), .ZN(n1582) );
  AOI221_X2 U910 ( .B1(ymem_data1[166]), .B2(n3292), .C1(ymem_data1[230]), 
        .C2(n3257), .A(n1583), .ZN(n1580) );
  OAI22_X2 U911 ( .A1(n3307), .A2(n332), .B1(n3284), .B2(n396), .ZN(n1583) );
  AOI221_X2 U913 ( .B1(ymem_data2[166]), .B2(n3271), .C1(ymem_data2[230]), 
        .C2(n849), .A(n1586), .ZN(n1585) );
  OAI22_X2 U914 ( .A1(n3266), .A2(n524), .B1(n3264), .B2(n588), .ZN(n1586) );
  AOI221_X2 U915 ( .B1(ymem_data1[38]), .B2(n3263), .C1(ymem_data1[102]), .C2(
        n854), .A(n1587), .ZN(n1584) );
  OAI22_X2 U916 ( .A1(n3259), .A2(n204), .B1(n3255), .B2(n268), .ZN(n1587) );
  AOI221_X2 U918 ( .B1(ymem_data1[38]), .B2(n3293), .C1(ymem_data2[230]), .C2(
        n3253), .A(n1590), .ZN(n1589) );
  OAI22_X2 U919 ( .A1(n3251), .A2(n332), .B1(n3249), .B2(n268), .ZN(n1590) );
  OAI22_X2 U922 ( .A1(n3240), .A2(n524), .B1(n99), .B2(n460), .ZN(n1592) );
  OAI221_X2 U923 ( .B1(n3248), .B2(n268), .C1(n3238), .C2(n332), .A(n1593), 
        .ZN(n1591) );
  OAI221_X2 U925 ( .B1(n1594), .B2(n3274), .C1(n3309), .C2(n19), .A(n1595), 
        .ZN(n2670) );
  AOI221_X2 U928 ( .B1(ymem_data2[167]), .B2(n3276), .C1(ymem_data2[231]), 
        .C2(n3297), .A(n1601), .ZN(n1600) );
  OAI22_X2 U929 ( .A1(n3305), .A2(n523), .B1(n3303), .B2(n587), .ZN(n1601) );
  AOI221_X2 U930 ( .B1(ymem_data1[167]), .B2(n3292), .C1(ymem_data1[231]), 
        .C2(n3257), .A(n1602), .ZN(n1599) );
  OAI22_X2 U931 ( .A1(n3307), .A2(n331), .B1(n3284), .B2(n395), .ZN(n1602) );
  AOI221_X2 U933 ( .B1(ymem_data2[167]), .B2(n3270), .C1(ymem_data2[231]), 
        .C2(n3268), .A(n1605), .ZN(n1604) );
  OAI22_X2 U934 ( .A1(n3266), .A2(n523), .B1(n3264), .B2(n587), .ZN(n1605) );
  AOI221_X2 U935 ( .B1(ymem_data1[39]), .B2(n3263), .C1(ymem_data1[103]), .C2(
        n3261), .A(n1606), .ZN(n1603) );
  OAI22_X2 U936 ( .A1(n3259), .A2(n203), .B1(n3255), .B2(n267), .ZN(n1606) );
  AOI221_X2 U938 ( .B1(ymem_data1[39]), .B2(n3293), .C1(ymem_data2[231]), .C2(
        n3253), .A(n1609), .ZN(n1608) );
  OAI22_X2 U939 ( .A1(n3251), .A2(n331), .B1(n3248), .B2(n267), .ZN(n1609) );
  OAI22_X2 U942 ( .A1(n3240), .A2(n523), .B1(n99), .B2(n459), .ZN(n1611) );
  OAI221_X2 U943 ( .B1(n863), .B2(n267), .C1(n3238), .C2(n331), .A(n1612), 
        .ZN(n1610) );
  OAI221_X2 U945 ( .B1(n1613), .B2(n3274), .C1(n3309), .C2(n18), .A(n1614), 
        .ZN(n2671) );
  AOI221_X2 U948 ( .B1(ymem_data2[168]), .B2(n3277), .C1(ymem_data2[232]), 
        .C2(n3296), .A(n1620), .ZN(n1619) );
  OAI22_X2 U949 ( .A1(n3305), .A2(n522), .B1(n3303), .B2(n586), .ZN(n1620) );
  AOI221_X2 U950 ( .B1(ymem_data1[168]), .B2(n3292), .C1(ymem_data1[232]), 
        .C2(n3257), .A(n1621), .ZN(n1618) );
  OAI22_X2 U951 ( .A1(n3307), .A2(n330), .B1(n3284), .B2(n394), .ZN(n1621) );
  AOI221_X2 U953 ( .B1(ymem_data2[168]), .B2(n3271), .C1(ymem_data2[232]), 
        .C2(n3268), .A(n1624), .ZN(n1623) );
  OAI22_X2 U954 ( .A1(n3266), .A2(n522), .B1(n3264), .B2(n586), .ZN(n1624) );
  AOI221_X2 U955 ( .B1(ymem_data1[40]), .B2(n3263), .C1(ymem_data1[104]), .C2(
        n854), .A(n1625), .ZN(n1622) );
  OAI22_X2 U956 ( .A1(n3259), .A2(n202), .B1(n3255), .B2(n266), .ZN(n1625) );
  AOI221_X2 U958 ( .B1(ymem_data1[40]), .B2(n3293), .C1(ymem_data2[232]), .C2(
        n3253), .A(n1628), .ZN(n1627) );
  OAI22_X2 U959 ( .A1(n3251), .A2(n330), .B1(n3249), .B2(n266), .ZN(n1628) );
  OAI22_X2 U962 ( .A1(n3240), .A2(n522), .B1(n99), .B2(n458), .ZN(n1630) );
  OAI221_X2 U963 ( .B1(n3249), .B2(n266), .C1(n3238), .C2(n330), .A(n1631), 
        .ZN(n1629) );
  OAI221_X2 U965 ( .B1(n1632), .B2(n3274), .C1(n3309), .C2(n17), .A(n1633), 
        .ZN(n2672) );
  AOI221_X2 U968 ( .B1(ymem_data2[169]), .B2(n3276), .C1(ymem_data2[233]), 
        .C2(n3297), .A(n1639), .ZN(n1638) );
  OAI22_X2 U969 ( .A1(n3305), .A2(n521), .B1(n3303), .B2(n585), .ZN(n1639) );
  AOI221_X2 U970 ( .B1(ymem_data1[169]), .B2(n3292), .C1(ymem_data1[233]), 
        .C2(n3257), .A(n1640), .ZN(n1637) );
  OAI22_X2 U971 ( .A1(n3307), .A2(n329), .B1(n778), .B2(n393), .ZN(n1640) );
  AOI221_X2 U973 ( .B1(ymem_data2[169]), .B2(n3270), .C1(ymem_data2[233]), 
        .C2(n3268), .A(n1643), .ZN(n1642) );
  OAI22_X2 U974 ( .A1(n3266), .A2(n521), .B1(n3264), .B2(n585), .ZN(n1643) );
  AOI221_X2 U975 ( .B1(ymem_data1[41]), .B2(n3263), .C1(ymem_data1[105]), .C2(
        n3261), .A(n1644), .ZN(n1641) );
  OAI22_X2 U976 ( .A1(n3259), .A2(n201), .B1(n3255), .B2(n265), .ZN(n1644) );
  AOI221_X2 U978 ( .B1(ymem_data1[41]), .B2(n3293), .C1(ymem_data2[233]), .C2(
        n3253), .A(n1647), .ZN(n1646) );
  OAI22_X2 U979 ( .A1(n3251), .A2(n329), .B1(n3248), .B2(n265), .ZN(n1647) );
  OAI22_X2 U982 ( .A1(n3240), .A2(n521), .B1(n99), .B2(n457), .ZN(n1649) );
  OAI221_X2 U983 ( .B1(n3248), .B2(n265), .C1(n3238), .C2(n329), .A(n1650), 
        .ZN(n1648) );
  OAI221_X2 U985 ( .B1(n1651), .B2(n3274), .C1(n3309), .C2(n16), .A(n1652), 
        .ZN(n2673) );
  AOI221_X2 U988 ( .B1(ymem_data2[170]), .B2(n3277), .C1(ymem_data2[234]), 
        .C2(n3296), .A(n1658), .ZN(n1657) );
  OAI22_X2 U989 ( .A1(n3305), .A2(n520), .B1(n3303), .B2(n584), .ZN(n1658) );
  AOI221_X2 U990 ( .B1(ymem_data1[170]), .B2(n3292), .C1(ymem_data1[234]), 
        .C2(n3257), .A(n1659), .ZN(n1656) );
  AOI221_X2 U993 ( .B1(ymem_data2[170]), .B2(n3271), .C1(ymem_data2[234]), 
        .C2(n3268), .A(n1662), .ZN(n1661) );
  OAI22_X2 U994 ( .A1(n3266), .A2(n520), .B1(n3264), .B2(n584), .ZN(n1662) );
  AOI221_X2 U995 ( .B1(ymem_data1[42]), .B2(n3263), .C1(ymem_data1[106]), .C2(
        n854), .A(n1663), .ZN(n1660) );
  OAI22_X2 U996 ( .A1(n3259), .A2(n200), .B1(n3255), .B2(n264), .ZN(n1663) );
  AOI221_X2 U998 ( .B1(ymem_data1[42]), .B2(n3293), .C1(ymem_data2[234]), .C2(
        n3253), .A(n1666), .ZN(n1665) );
  OAI22_X2 U999 ( .A1(n3251), .A2(n328), .B1(n3249), .B2(n264), .ZN(n1666) );
  OAI22_X2 U1002 ( .A1(n3240), .A2(n520), .B1(n99), .B2(n456), .ZN(n1668) );
  OAI221_X2 U1003 ( .B1(n3248), .B2(n264), .C1(n3238), .C2(n328), .A(n1669), 
        .ZN(n1667) );
  OAI221_X2 U1005 ( .B1(n1670), .B2(n3274), .C1(n3309), .C2(n15), .A(n1671), 
        .ZN(n2674) );
  AOI221_X2 U1008 ( .B1(ymem_data2[171]), .B2(n3276), .C1(ymem_data2[235]), 
        .C2(n3296), .A(n1677), .ZN(n1676) );
  OAI22_X2 U1009 ( .A1(n3305), .A2(n519), .B1(n3303), .B2(n583), .ZN(n1677) );
  AOI221_X2 U1010 ( .B1(ymem_data1[171]), .B2(n3292), .C1(ymem_data1[235]), 
        .C2(n3258), .A(n1678), .ZN(n1675) );
  AOI221_X2 U1013 ( .B1(ymem_data2[171]), .B2(n3270), .C1(ymem_data2[235]), 
        .C2(n3268), .A(n1681), .ZN(n1680) );
  OAI22_X2 U1014 ( .A1(n3266), .A2(n519), .B1(n3264), .B2(n583), .ZN(n1681) );
  AOI221_X2 U1015 ( .B1(ymem_data1[43]), .B2(n3263), .C1(ymem_data1[107]), 
        .C2(n3261), .A(n1682), .ZN(n1679) );
  OAI22_X2 U1016 ( .A1(n856), .A2(n199), .B1(n3255), .B2(n263), .ZN(n1682) );
  AOI221_X2 U1018 ( .B1(ymem_data1[43]), .B2(n3293), .C1(ymem_data2[235]), 
        .C2(n3253), .A(n1685), .ZN(n1684) );
  OAI22_X2 U1019 ( .A1(n3251), .A2(n327), .B1(n3248), .B2(n263), .ZN(n1685) );
  OAI22_X2 U1022 ( .A1(n3240), .A2(n519), .B1(n99), .B2(n455), .ZN(n1687) );
  OAI221_X2 U1023 ( .B1(n3248), .B2(n263), .C1(n3238), .C2(n327), .A(n1688), 
        .ZN(n1686) );
  OAI221_X2 U1025 ( .B1(n1689), .B2(n3274), .C1(n3309), .C2(n14), .A(n1690), 
        .ZN(n2675) );
  AOI221_X2 U1028 ( .B1(ymem_data2[172]), .B2(n3277), .C1(ymem_data2[236]), 
        .C2(n3297), .A(n1696), .ZN(n1695) );
  OAI22_X2 U1029 ( .A1(n3305), .A2(n518), .B1(n3303), .B2(n582), .ZN(n1696) );
  AOI221_X2 U1030 ( .B1(ymem_data1[172]), .B2(n110), .C1(ymem_data1[236]), 
        .C2(n3257), .A(n1697), .ZN(n1694) );
  AOI221_X2 U1033 ( .B1(ymem_data2[172]), .B2(n3271), .C1(ymem_data2[236]), 
        .C2(n3268), .A(n1700), .ZN(n1699) );
  OAI22_X2 U1034 ( .A1(n3266), .A2(n518), .B1(n3264), .B2(n582), .ZN(n1700) );
  AOI221_X2 U1035 ( .B1(ymem_data1[44]), .B2(n3263), .C1(ymem_data1[108]), 
        .C2(n3261), .A(n1701), .ZN(n1698) );
  OAI22_X2 U1036 ( .A1(n3259), .A2(n198), .B1(n3255), .B2(n262), .ZN(n1701) );
  AOI221_X2 U1038 ( .B1(ymem_data1[44]), .B2(n3293), .C1(ymem_data2[236]), 
        .C2(n3253), .A(n1704), .ZN(n1703) );
  OAI22_X2 U1039 ( .A1(n3251), .A2(n326), .B1(n3249), .B2(n262), .ZN(n1704) );
  OAI22_X2 U1042 ( .A1(n3240), .A2(n518), .B1(n99), .B2(n454), .ZN(n1706) );
  OAI221_X2 U1045 ( .B1(n1708), .B2(n3274), .C1(n3309), .C2(n13), .A(n1709), 
        .ZN(n2676) );
  AOI221_X2 U1048 ( .B1(ymem_data2[173]), .B2(n3276), .C1(ymem_data2[237]), 
        .C2(n3297), .A(n1715), .ZN(n1714) );
  OAI22_X2 U1049 ( .A1(n3305), .A2(n517), .B1(n3303), .B2(n581), .ZN(n1715) );
  AOI221_X2 U1050 ( .B1(ymem_data1[173]), .B2(n110), .C1(ymem_data1[237]), 
        .C2(n3257), .A(n1716), .ZN(n1713) );
  OAI22_X2 U1051 ( .A1(n3307), .A2(n325), .B1(n3284), .B2(n389), .ZN(n1716) );
  AOI221_X2 U1053 ( .B1(ymem_data2[173]), .B2(n3270), .C1(ymem_data2[237]), 
        .C2(n3268), .A(n1719), .ZN(n1718) );
  OAI22_X2 U1054 ( .A1(n3266), .A2(n517), .B1(n3264), .B2(n581), .ZN(n1719) );
  AOI221_X2 U1055 ( .B1(ymem_data1[45]), .B2(n3263), .C1(ymem_data1[109]), 
        .C2(n3261), .A(n1720), .ZN(n1717) );
  OAI22_X2 U1056 ( .A1(n3259), .A2(n197), .B1(n3255), .B2(n261), .ZN(n1720) );
  AOI221_X2 U1058 ( .B1(ymem_data1[45]), .B2(n3293), .C1(ymem_data2[237]), 
        .C2(n3253), .A(n1723), .ZN(n1722) );
  OAI22_X2 U1059 ( .A1(n3251), .A2(n325), .B1(n3248), .B2(n261), .ZN(n1723) );
  OAI22_X2 U1062 ( .A1(n3240), .A2(n517), .B1(n99), .B2(n453), .ZN(n1725) );
  OAI221_X2 U1063 ( .B1(n3248), .B2(n261), .C1(n3238), .C2(n325), .A(n1726), 
        .ZN(n1724) );
  OAI221_X2 U1065 ( .B1(n1727), .B2(n3274), .C1(n3309), .C2(n12), .A(n1728), 
        .ZN(n2677) );
  AOI221_X2 U1068 ( .B1(ymem_data2[174]), .B2(n3277), .C1(ymem_data2[238]), 
        .C2(n3296), .A(n1734), .ZN(n1733) );
  OAI22_X2 U1069 ( .A1(n3305), .A2(n516), .B1(n3303), .B2(n580), .ZN(n1734) );
  AOI221_X2 U1070 ( .B1(ymem_data1[174]), .B2(n110), .C1(ymem_data1[238]), 
        .C2(n3257), .A(n1735), .ZN(n1732) );
  OAI22_X2 U1071 ( .A1(n3307), .A2(n324), .B1(n3284), .B2(n388), .ZN(n1735) );
  AOI221_X2 U1073 ( .B1(ymem_data2[174]), .B2(n3271), .C1(ymem_data2[238]), 
        .C2(n3268), .A(n1738), .ZN(n1737) );
  OAI22_X2 U1074 ( .A1(n3266), .A2(n516), .B1(n3264), .B2(n580), .ZN(n1738) );
  AOI221_X2 U1075 ( .B1(ymem_data1[46]), .B2(n3263), .C1(ymem_data1[110]), 
        .C2(n3261), .A(n1739), .ZN(n1736) );
  OAI22_X2 U1076 ( .A1(n3259), .A2(n196), .B1(n3255), .B2(n260), .ZN(n1739) );
  AOI221_X2 U1078 ( .B1(ymem_data1[46]), .B2(n3293), .C1(ymem_data2[238]), 
        .C2(n3253), .A(n1742), .ZN(n1741) );
  OAI22_X2 U1079 ( .A1(n3251), .A2(n324), .B1(n3248), .B2(n260), .ZN(n1742) );
  OAI22_X2 U1082 ( .A1(n3240), .A2(n516), .B1(n99), .B2(n452), .ZN(n1744) );
  OAI221_X2 U1085 ( .B1(n1746), .B2(n3274), .C1(n3309), .C2(n11), .A(n1747), 
        .ZN(n2678) );
  AOI221_X2 U1089 ( .B1(ymem_data2[175]), .B2(n3276), .C1(ymem_data2[239]), 
        .C2(n3297), .A(n1754), .ZN(n1752) );
  OAI22_X2 U1090 ( .A1(n3305), .A2(n515), .B1(n3303), .B2(n579), .ZN(n1754) );
  NAND2_X2 U1093 ( .A1(n712), .A2(n3259), .ZN(n723) );
  AOI221_X2 U1095 ( .B1(ymem_data1[175]), .B2(n110), .C1(ymem_data1[239]), 
        .C2(n3257), .A(n1755), .ZN(n1751) );
  OAI22_X2 U1096 ( .A1(n3307), .A2(n323), .B1(n3284), .B2(n387), .ZN(n1755) );
  NAND2_X2 U1097 ( .A1(n699), .A2(n3259), .ZN(n778) );
  NAND2_X2 U1099 ( .A1(n111), .A2(n3259), .ZN(n815) );
  AOI221_X2 U1102 ( .B1(ymem_data2[175]), .B2(n3270), .C1(ymem_data2[239]), 
        .C2(n3268), .A(n1758), .ZN(n1757) );
  OAI22_X2 U1103 ( .A1(n3266), .A2(n515), .B1(n3264), .B2(n579), .ZN(n1758) );
  AOI221_X2 U1104 ( .B1(ymem_data1[47]), .B2(n3263), .C1(ymem_data1[111]), 
        .C2(n3261), .A(n1759), .ZN(n1756) );
  OAI22_X2 U1105 ( .A1(n3259), .A2(n195), .B1(n3255), .B2(n259), .ZN(n1759) );
  AOI221_X2 U1107 ( .B1(ymem_data1[47]), .B2(n3293), .C1(ymem_data2[239]), 
        .C2(n3253), .A(n1762), .ZN(n1761) );
  OAI22_X2 U1108 ( .A1(n3251), .A2(n323), .B1(n3249), .B2(n259), .ZN(n1762) );
  OAI221_X2 U1110 ( .B1(n697), .B2(n711), .C1(n3203), .C2(n707), .A(n1763), 
        .ZN(n860) );
  NOR2_X2 U1112 ( .A1(n707), .A2(n109), .ZN(n712) );
  OAI221_X2 U1115 ( .B1(n701), .B2(n796), .C1(n697), .C2(n709), .A(n1765), 
        .ZN(n865) );
  NAND2_X2 U1117 ( .A1(n749), .A2(n1766), .ZN(n706) );
  NAND2_X2 U1118 ( .A1(n799), .A2(n698), .ZN(n709) );
  OAI221_X2 U1119 ( .B1(n701), .B2(n102), .C1(n697), .C2(n710), .A(n1767), 
        .ZN(n864) );
  OAI221_X2 U1120 ( .B1(n701), .B2(n1769), .C1(n697), .C2(n708), .A(n1770), 
        .ZN(n1768) );
  NAND2_X2 U1122 ( .A1(n94), .A2(n1771), .ZN(n708) );
  NOR2_X2 U1125 ( .A1(n9), .A2(n131), .ZN(n828) );
  OAI22_X2 U1127 ( .A1(n3240), .A2(n515), .B1(n99), .B2(n451), .ZN(n1774) );
  OAI221_X2 U1128 ( .B1(n734), .B2(n747), .C1(n739), .C2(n102), .A(n1767), 
        .ZN(n1775) );
  NAND2_X2 U1130 ( .A1(n745), .A2(n698), .ZN(n814) );
  NOR2_X2 U1131 ( .A1(n747), .A2(n132), .ZN(n745) );
  NAND2_X2 U1132 ( .A1(n1776), .A2(n735), .ZN(n747) );
  AOI221_X2 U1133 ( .B1(n120), .B2(n799), .C1(n115), .C2(n749), .A(n1777), 
        .ZN(n869) );
  OAI22_X2 U1134 ( .A1(n744), .A2(n3203), .B1(n96), .B2(n695), .ZN(n1777) );
  NOR2_X2 U1135 ( .A1(n744), .A2(n109), .ZN(n751) );
  NAND2_X2 U1136 ( .A1(n799), .A2(n728), .ZN(n744) );
  NOR2_X2 U1137 ( .A1(n796), .A2(n111), .ZN(n749) );
  NAND2_X2 U1138 ( .A1(n109), .A2(n1778), .ZN(n796) );
  OAI221_X2 U1139 ( .B1(n3248), .B2(n259), .C1(n3238), .C2(n323), .A(n1779), 
        .ZN(n1773) );
  AOI221_X2 U1141 ( .B1(n146), .B2(n750), .C1(n115), .C2(n105), .A(n1781), 
        .ZN(n1780) );
  OAI22_X2 U1142 ( .A1(n707), .A2(n3203), .B1(n825), .B2(n739), .ZN(n1781) );
  NAND2_X2 U1143 ( .A1(n105), .A2(n1766), .ZN(n707) );
  NOR3_X2 U1144 ( .A1(n107), .A2(n109), .A3(n792), .ZN(n750) );
  NAND2_X2 U1145 ( .A1(n132), .A2(n735), .ZN(n792) );
  NOR3_X2 U1147 ( .A1(n107), .A2(n111), .A3(n698), .ZN(n736) );
  NAND2_X2 U1149 ( .A1(n107), .A2(n735), .ZN(n748) );
  NAND2_X2 U1150 ( .A1(n111), .A2(n146), .ZN(n863) );
  OAI221_X2 U1151 ( .B1(n739), .B2(n1783), .C1(n734), .C2(n746), .A(n1784), 
        .ZN(n866) );
  NOR2_X2 U1153 ( .A1(n93), .A2(n118), .ZN(n752) );
  NOR2_X2 U1154 ( .A1(n746), .A2(n132), .ZN(n784) );
  NAND2_X2 U1155 ( .A1(n91), .A2(n728), .ZN(n743) );
  NAND2_X2 U1156 ( .A1(n94), .A2(n735), .ZN(n746) );
  NAND3_X2 U1157 ( .A1(n1778), .A2(n698), .A3(n95), .ZN(n1769) );
  NAND3_X2 U1158 ( .A1(n1778), .A2(n1771), .A3(n95), .ZN(n1783) );
  AND4_X2 U1160 ( .A1(n829), .A2(n717), .A3(n634), .A4(n1786), .ZN(n1785) );
  NOR4_X2 U1163 ( .A1(n780), .A2(n804), .A3(n813), .A4(n4), .ZN(n714) );
  NOR4_X2 U1164 ( .A1(n5), .A2(n805), .A3(n812), .A4(n727), .ZN(n724) );
  AOI221_X2 U1166 ( .B1(yMemDataReadyNextCycle), .B2(n3215), .C1(n3287), .C2(
        n1792), .A(n130), .ZN(n1790) );
  NOR4_X2 U1168 ( .A1(n1795), .A2(n1796), .A3(n3202), .A4(n3291), .ZN(n1793)
         );
  AND3_X2 U1169 ( .A1(n1798), .A2(n152), .A3(filt_EN), .ZN(n1796) );
  NAND2_X2 U1171 ( .A1(n3), .A2(exModDone), .ZN(n1792) );
  AOI221_X2 U1174 ( .B1(ymem_data1[201]), .B2(n3282), .C1(ymem_data1[137]), 
        .C2(n3280), .A(n1803), .ZN(n1801) );
  AOI221_X2 U1176 ( .B1(n3235), .B2(ymem_data2[201]), .C1(n3232), .C2(
        ymem_data1[9]), .A(n1808), .ZN(n1805) );
  AOI221_X2 U1178 ( .B1(n3225), .B2(ymem_data1[201]), .C1(n3236), .C2(
        U72_DATA1_9), .A(n1813), .ZN(n1804) );
  OAI22_X2 U1179 ( .A1(n297), .A2(n3198), .B1(n361), .B2(n1815), .ZN(n1813) );
  AOI221_X2 U1182 ( .B1(ymem_data1[200]), .B2(n3282), .C1(ymem_data1[136]), 
        .C2(n3280), .A(n1818), .ZN(n1816) );
  AOI221_X2 U1184 ( .B1(n3234), .B2(ymem_data2[200]), .C1(n3232), .C2(
        ymem_data1[8]), .A(n1821), .ZN(n1820) );
  AOI221_X2 U1186 ( .B1(n3224), .B2(ymem_data1[200]), .C1(n3236), .C2(
        U72_DATA1_8), .A(n1822), .ZN(n1819) );
  OAI22_X2 U1187 ( .A1(n298), .A2(n3198), .B1(n362), .B2(n1815), .ZN(n1822) );
  AOI221_X2 U1190 ( .B1(ymem_data1[199]), .B2(n3282), .C1(ymem_data1[135]), 
        .C2(n3280), .A(n1825), .ZN(n1823) );
  AOI221_X2 U1192 ( .B1(n3235), .B2(ymem_data2[199]), .C1(n1807), .C2(
        ymem_data1[7]), .A(n1828), .ZN(n1827) );
  AOI221_X2 U1194 ( .B1(n3225), .B2(ymem_data1[199]), .C1(n3236), .C2(
        U72_DATA1_7), .A(n1829), .ZN(n1826) );
  OAI22_X2 U1195 ( .A1(n299), .A2(n3198), .B1(n363), .B2(n1815), .ZN(n1829) );
  AOI221_X2 U1198 ( .B1(ymem_data1[198]), .B2(n3282), .C1(ymem_data1[134]), 
        .C2(n3280), .A(n1832), .ZN(n1830) );
  AOI221_X2 U1200 ( .B1(n3234), .B2(ymem_data2[198]), .C1(n1807), .C2(
        ymem_data1[6]), .A(n1835), .ZN(n1834) );
  AOI221_X2 U1202 ( .B1(n3224), .B2(ymem_data1[198]), .C1(n3236), .C2(
        U72_DATA1_6), .A(n1836), .ZN(n1833) );
  OAI22_X2 U1203 ( .A1(n300), .A2(n3198), .B1(n364), .B2(n1815), .ZN(n1836) );
  AOI221_X2 U1206 ( .B1(ymem_data1[197]), .B2(n3282), .C1(ymem_data1[133]), 
        .C2(n3280), .A(n1839), .ZN(n1837) );
  AOI221_X2 U1208 ( .B1(n3235), .B2(ymem_data2[197]), .C1(n1807), .C2(
        ymem_data1[5]), .A(n1842), .ZN(n1841) );
  AOI221_X2 U1210 ( .B1(n3224), .B2(ymem_data1[197]), .C1(n3236), .C2(
        U72_DATA1_5), .A(n1843), .ZN(n1840) );
  OAI22_X2 U1211 ( .A1(n301), .A2(n3198), .B1(n365), .B2(n1815), .ZN(n1843) );
  AOI221_X2 U1214 ( .B1(ymem_data1[239]), .B2(n3282), .C1(ymem_data1[175]), 
        .C2(n3280), .A(n1846), .ZN(n1844) );
  AOI221_X2 U1216 ( .B1(n3234), .B2(ymem_data2[239]), .C1(n1807), .C2(
        ymem_data1[47]), .A(n1849), .ZN(n1848) );
  AOI221_X2 U1218 ( .B1(n3225), .B2(ymem_data1[239]), .C1(n3236), .C2(
        U72_DATA1_47), .A(n1850), .ZN(n1847) );
  OAI22_X2 U1219 ( .A1(n259), .A2(n3198), .B1(n323), .B2(n1815), .ZN(n1850) );
  AOI221_X2 U1222 ( .B1(ymem_data1[238]), .B2(n3282), .C1(ymem_data1[174]), 
        .C2(n3280), .A(n1853), .ZN(n1851) );
  AOI221_X2 U1224 ( .B1(n3234), .B2(ymem_data2[238]), .C1(n1807), .C2(
        ymem_data1[46]), .A(n1856), .ZN(n1855) );
  AOI221_X2 U1226 ( .B1(n3225), .B2(ymem_data1[238]), .C1(n3236), .C2(
        U72_DATA1_46), .A(n1857), .ZN(n1854) );
  OAI22_X2 U1227 ( .A1(n260), .A2(n3198), .B1(n324), .B2(n1815), .ZN(n1857) );
  AOI221_X2 U1230 ( .B1(ymem_data1[237]), .B2(n3282), .C1(ymem_data1[173]), 
        .C2(n3280), .A(n1860), .ZN(n1858) );
  AOI221_X2 U1232 ( .B1(n3235), .B2(ymem_data2[237]), .C1(n1807), .C2(
        ymem_data1[45]), .A(n1863), .ZN(n1862) );
  AOI221_X2 U1234 ( .B1(n3224), .B2(ymem_data1[237]), .C1(n3236), .C2(
        U72_DATA1_45), .A(n1864), .ZN(n1861) );
  OAI22_X2 U1235 ( .A1(n261), .A2(n3198), .B1(n325), .B2(n1815), .ZN(n1864) );
  AOI221_X2 U1238 ( .B1(ymem_data1[236]), .B2(n3282), .C1(ymem_data1[172]), 
        .C2(n3280), .A(n1867), .ZN(n1865) );
  AOI221_X2 U1240 ( .B1(n3234), .B2(ymem_data2[236]), .C1(n1807), .C2(
        ymem_data1[44]), .A(n1870), .ZN(n1869) );
  AOI221_X2 U1242 ( .B1(n3225), .B2(ymem_data1[236]), .C1(n3236), .C2(
        U72_DATA1_44), .A(n1871), .ZN(n1868) );
  OAI22_X2 U1243 ( .A1(n262), .A2(n3198), .B1(n326), .B2(n3223), .ZN(n1871) );
  AOI221_X2 U1246 ( .B1(ymem_data1[235]), .B2(n3282), .C1(ymem_data1[171]), 
        .C2(n3280), .A(n1874), .ZN(n1872) );
  AOI221_X2 U1248 ( .B1(n3235), .B2(ymem_data2[235]), .C1(n1807), .C2(
        ymem_data1[43]), .A(n1877), .ZN(n1876) );
  AOI221_X2 U1250 ( .B1(n3224), .B2(ymem_data1[235]), .C1(n3236), .C2(
        U72_DATA1_43), .A(n1878), .ZN(n1875) );
  OAI22_X2 U1251 ( .A1(n263), .A2(n3198), .B1(n327), .B2(n3223), .ZN(n1878) );
  AOI221_X2 U1254 ( .B1(ymem_data1[234]), .B2(n3282), .C1(ymem_data1[170]), 
        .C2(n3280), .A(n1881), .ZN(n1879) );
  AOI221_X2 U1256 ( .B1(n3235), .B2(ymem_data2[234]), .C1(n1807), .C2(
        ymem_data1[42]), .A(n1884), .ZN(n1883) );
  AOI221_X2 U1258 ( .B1(n3225), .B2(ymem_data1[234]), .C1(n3236), .C2(
        U72_DATA1_42), .A(n1885), .ZN(n1882) );
  OAI22_X2 U1259 ( .A1(n264), .A2(n3198), .B1(n328), .B2(n3223), .ZN(n1885) );
  AOI221_X2 U1262 ( .B1(ymem_data1[233]), .B2(n3282), .C1(ymem_data1[169]), 
        .C2(n3280), .A(n1888), .ZN(n1886) );
  AOI221_X2 U1264 ( .B1(n3235), .B2(ymem_data2[233]), .C1(n1807), .C2(
        ymem_data1[41]), .A(n1891), .ZN(n1890) );
  AOI221_X2 U1266 ( .B1(n3224), .B2(ymem_data1[233]), .C1(n3236), .C2(
        U72_DATA1_41), .A(n1892), .ZN(n1889) );
  OAI22_X2 U1267 ( .A1(n265), .A2(n3198), .B1(n329), .B2(n3223), .ZN(n1892) );
  AOI221_X2 U1270 ( .B1(ymem_data1[232]), .B2(n3282), .C1(ymem_data1[168]), 
        .C2(n3280), .A(n1895), .ZN(n1893) );
  AOI221_X2 U1272 ( .B1(n3235), .B2(ymem_data2[232]), .C1(n1807), .C2(
        ymem_data1[40]), .A(n1898), .ZN(n1897) );
  AOI221_X2 U1274 ( .B1(n3225), .B2(ymem_data1[232]), .C1(n3236), .C2(
        U72_DATA1_40), .A(n1899), .ZN(n1896) );
  OAI22_X2 U1275 ( .A1(n266), .A2(n3198), .B1(n330), .B2(n3223), .ZN(n1899) );
  AOI221_X2 U1278 ( .B1(ymem_data1[196]), .B2(n3282), .C1(ymem_data1[132]), 
        .C2(n3280), .A(n1902), .ZN(n1900) );
  AOI221_X2 U1280 ( .B1(n3235), .B2(ymem_data2[196]), .C1(n1807), .C2(
        ymem_data1[4]), .A(n1905), .ZN(n1904) );
  AOI221_X2 U1282 ( .B1(n3224), .B2(ymem_data1[196]), .C1(n3236), .C2(
        U72_DATA1_4), .A(n1906), .ZN(n1903) );
  OAI22_X2 U1283 ( .A1(n302), .A2(n3198), .B1(n366), .B2(n3223), .ZN(n1906) );
  AOI221_X2 U1286 ( .B1(ymem_data1[231]), .B2(n3282), .C1(ymem_data1[167]), 
        .C2(n3280), .A(n1909), .ZN(n1907) );
  AOI221_X2 U1288 ( .B1(n3235), .B2(ymem_data2[231]), .C1(n3232), .C2(
        ymem_data1[39]), .A(n1912), .ZN(n1911) );
  AOI221_X2 U1290 ( .B1(n3225), .B2(ymem_data1[231]), .C1(n3236), .C2(
        U72_DATA1_39), .A(n1913), .ZN(n1910) );
  OAI22_X2 U1291 ( .A1(n267), .A2(n3198), .B1(n331), .B2(n3223), .ZN(n1913) );
  AOI221_X2 U1294 ( .B1(ymem_data1[230]), .B2(n3282), .C1(ymem_data1[166]), 
        .C2(n3280), .A(n1916), .ZN(n1914) );
  AOI221_X2 U1296 ( .B1(n3235), .B2(ymem_data2[230]), .C1(n3232), .C2(
        ymem_data1[38]), .A(n1919), .ZN(n1918) );
  AOI221_X2 U1298 ( .B1(n3224), .B2(ymem_data1[230]), .C1(n3236), .C2(
        U72_DATA1_38), .A(n1920), .ZN(n1917) );
  OAI22_X2 U1299 ( .A1(n268), .A2(n3198), .B1(n332), .B2(n3223), .ZN(n1920) );
  AOI221_X2 U1302 ( .B1(ymem_data1[229]), .B2(n3282), .C1(ymem_data1[165]), 
        .C2(n3280), .A(n1923), .ZN(n1921) );
  AOI221_X2 U1304 ( .B1(n3235), .B2(ymem_data2[229]), .C1(n3232), .C2(
        ymem_data1[37]), .A(n1926), .ZN(n1925) );
  AOI221_X2 U1306 ( .B1(n3225), .B2(ymem_data1[229]), .C1(n3236), .C2(
        U72_DATA1_37), .A(n1927), .ZN(n1924) );
  OAI22_X2 U1307 ( .A1(n269), .A2(n3198), .B1(n333), .B2(n3223), .ZN(n1927) );
  AOI221_X2 U1310 ( .B1(ymem_data1[228]), .B2(n3282), .C1(ymem_data1[164]), 
        .C2(n3280), .A(n1930), .ZN(n1928) );
  AOI221_X2 U1312 ( .B1(n3235), .B2(ymem_data2[228]), .C1(n3232), .C2(
        ymem_data1[36]), .A(n1933), .ZN(n1932) );
  AOI221_X2 U1314 ( .B1(n3224), .B2(ymem_data1[228]), .C1(n3236), .C2(
        U72_DATA1_36), .A(n1934), .ZN(n1931) );
  OAI22_X2 U1315 ( .A1(n270), .A2(n3198), .B1(n334), .B2(n3223), .ZN(n1934) );
  AOI221_X2 U1318 ( .B1(ymem_data1[227]), .B2(n3282), .C1(ymem_data1[163]), 
        .C2(n782), .A(n1937), .ZN(n1935) );
  AOI221_X2 U1320 ( .B1(n3235), .B2(ymem_data2[227]), .C1(n3232), .C2(
        ymem_data1[35]), .A(n1940), .ZN(n1939) );
  AOI221_X2 U1322 ( .B1(n3225), .B2(ymem_data1[227]), .C1(n3236), .C2(
        U72_DATA1_35), .A(n1941), .ZN(n1938) );
  OAI22_X2 U1323 ( .A1(n271), .A2(n3198), .B1(n335), .B2(n3223), .ZN(n1941) );
  AOI221_X2 U1326 ( .B1(ymem_data1[226]), .B2(n3282), .C1(ymem_data1[162]), 
        .C2(n782), .A(n1944), .ZN(n1942) );
  AOI221_X2 U1328 ( .B1(n3235), .B2(ymem_data2[226]), .C1(n3232), .C2(
        ymem_data1[34]), .A(n1947), .ZN(n1946) );
  AOI221_X2 U1330 ( .B1(n3224), .B2(ymem_data1[226]), .C1(n3236), .C2(
        U72_DATA1_34), .A(n1948), .ZN(n1945) );
  OAI22_X2 U1331 ( .A1(n272), .A2(n3198), .B1(n336), .B2(n3223), .ZN(n1948) );
  AOI221_X2 U1334 ( .B1(ymem_data1[225]), .B2(n3282), .C1(ymem_data1[161]), 
        .C2(n782), .A(n1951), .ZN(n1949) );
  AOI221_X2 U1336 ( .B1(n3235), .B2(ymem_data2[225]), .C1(n3232), .C2(
        ymem_data1[33]), .A(n1954), .ZN(n1953) );
  AOI221_X2 U1338 ( .B1(n3225), .B2(ymem_data1[225]), .C1(n3237), .C2(
        U72_DATA1_33), .A(n1955), .ZN(n1952) );
  OAI22_X2 U1339 ( .A1(n273), .A2(n3198), .B1(n337), .B2(n3223), .ZN(n1955) );
  AOI221_X2 U1342 ( .B1(ymem_data1[224]), .B2(n3282), .C1(ymem_data1[160]), 
        .C2(n3280), .A(n1958), .ZN(n1956) );
  AOI221_X2 U1344 ( .B1(n3235), .B2(ymem_data2[224]), .C1(n3232), .C2(
        ymem_data1[32]), .A(n1961), .ZN(n1960) );
  AOI221_X2 U1346 ( .B1(n3224), .B2(ymem_data1[224]), .C1(n3237), .C2(
        U72_DATA1_32), .A(n1962), .ZN(n1959) );
  OAI22_X2 U1347 ( .A1(n274), .A2(n3198), .B1(n338), .B2(n3223), .ZN(n1962) );
  AOI221_X2 U1350 ( .B1(ymem_data1[223]), .B2(n3283), .C1(ymem_data1[159]), 
        .C2(n3280), .A(n1965), .ZN(n1963) );
  AOI221_X2 U1352 ( .B1(n3234), .B2(ymem_data2[223]), .C1(n3232), .C2(
        ymem_data1[31]), .A(n1968), .ZN(n1967) );
  AOI221_X2 U1354 ( .B1(n3225), .B2(ymem_data1[223]), .C1(n3237), .C2(
        U72_DATA1_31), .A(n1969), .ZN(n1966) );
  OAI22_X2 U1355 ( .A1(n275), .A2(n3198), .B1(n339), .B2(n3223), .ZN(n1969) );
  AOI221_X2 U1358 ( .B1(ymem_data1[222]), .B2(n3283), .C1(ymem_data1[158]), 
        .C2(n3280), .A(n1972), .ZN(n1970) );
  AOI221_X2 U1360 ( .B1(n3234), .B2(ymem_data2[222]), .C1(n3232), .C2(
        ymem_data1[30]), .A(n1975), .ZN(n1974) );
  AOI221_X2 U1362 ( .B1(n3225), .B2(ymem_data1[222]), .C1(n3237), .C2(
        U72_DATA1_30), .A(n1976), .ZN(n1973) );
  OAI22_X2 U1363 ( .A1(n276), .A2(n3198), .B1(n340), .B2(n3223), .ZN(n1976) );
  AOI221_X2 U1366 ( .B1(ymem_data1[195]), .B2(n3283), .C1(ymem_data1[131]), 
        .C2(n3280), .A(n1979), .ZN(n1977) );
  AOI221_X2 U1368 ( .B1(n3234), .B2(ymem_data2[195]), .C1(n3232), .C2(
        ymem_data1[3]), .A(n1982), .ZN(n1981) );
  AOI221_X2 U1370 ( .B1(n3225), .B2(ymem_data1[195]), .C1(n3237), .C2(
        U72_DATA1_3), .A(n1983), .ZN(n1980) );
  OAI22_X2 U1371 ( .A1(n303), .A2(n3198), .B1(n367), .B2(n3223), .ZN(n1983) );
  AOI221_X2 U1374 ( .B1(ymem_data1[221]), .B2(n3283), .C1(ymem_data1[157]), 
        .C2(n782), .A(n1986), .ZN(n1984) );
  AOI221_X2 U1376 ( .B1(n3234), .B2(ymem_data2[221]), .C1(n3232), .C2(
        ymem_data1[29]), .A(n1989), .ZN(n1988) );
  AOI221_X2 U1378 ( .B1(n3225), .B2(ymem_data1[221]), .C1(n3237), .C2(
        U72_DATA1_29), .A(n1990), .ZN(n1987) );
  OAI22_X2 U1379 ( .A1(n277), .A2(n3198), .B1(n341), .B2(n1815), .ZN(n1990) );
  AOI221_X2 U1382 ( .B1(ymem_data1[220]), .B2(n3283), .C1(ymem_data1[156]), 
        .C2(n782), .A(n1993), .ZN(n1991) );
  AOI221_X2 U1384 ( .B1(n3234), .B2(ymem_data2[220]), .C1(n3232), .C2(
        ymem_data1[28]), .A(n1996), .ZN(n1995) );
  AOI221_X2 U1386 ( .B1(n3225), .B2(ymem_data1[220]), .C1(n3237), .C2(
        U72_DATA1_28), .A(n1997), .ZN(n1994) );
  OAI22_X2 U1387 ( .A1(n278), .A2(n3198), .B1(n342), .B2(n1815), .ZN(n1997) );
  AOI221_X2 U1392 ( .B1(n3234), .B2(ymem_data2[219]), .C1(n3232), .C2(
        ymem_data1[27]), .A(n2003), .ZN(n2002) );
  AOI221_X2 U1394 ( .B1(n3225), .B2(ymem_data1[219]), .C1(n3237), .C2(
        U72_DATA1_27), .A(n2004), .ZN(n2001) );
  OAI22_X2 U1395 ( .A1(n279), .A2(n3198), .B1(n343), .B2(n1815), .ZN(n2004) );
  AOI221_X2 U1398 ( .B1(ymem_data1[218]), .B2(n3283), .C1(ymem_data1[154]), 
        .C2(n782), .A(n2007), .ZN(n2005) );
  AOI221_X2 U1400 ( .B1(n3234), .B2(ymem_data2[218]), .C1(n3232), .C2(
        ymem_data1[26]), .A(n2010), .ZN(n2009) );
  AOI221_X2 U1402 ( .B1(n3225), .B2(ymem_data1[218]), .C1(n3237), .C2(
        U72_DATA1_26), .A(n2011), .ZN(n2008) );
  OAI22_X2 U1403 ( .A1(n280), .A2(n3198), .B1(n344), .B2(n3223), .ZN(n2011) );
  AOI221_X2 U1406 ( .B1(ymem_data1[217]), .B2(n3283), .C1(ymem_data1[153]), 
        .C2(n782), .A(n2014), .ZN(n2012) );
  AOI221_X2 U1408 ( .B1(n3234), .B2(ymem_data2[217]), .C1(n3232), .C2(
        ymem_data1[25]), .A(n2017), .ZN(n2016) );
  AOI221_X2 U1410 ( .B1(n3225), .B2(ymem_data1[217]), .C1(n3237), .C2(
        U72_DATA1_25), .A(n2018), .ZN(n2015) );
  OAI22_X2 U1411 ( .A1(n281), .A2(n3198), .B1(n345), .B2(n3223), .ZN(n2018) );
  AOI221_X2 U1414 ( .B1(ymem_data1[216]), .B2(n3283), .C1(ymem_data1[152]), 
        .C2(n782), .A(n2021), .ZN(n2019) );
  AOI221_X2 U1416 ( .B1(n3234), .B2(ymem_data2[216]), .C1(n3232), .C2(
        ymem_data1[24]), .A(n2024), .ZN(n2023) );
  AOI221_X2 U1418 ( .B1(n3225), .B2(ymem_data1[216]), .C1(n3237), .C2(
        U72_DATA1_24), .A(n2025), .ZN(n2022) );
  OAI22_X2 U1419 ( .A1(n282), .A2(n3198), .B1(n346), .B2(n1815), .ZN(n2025) );
  AOI221_X2 U1422 ( .B1(ymem_data1[215]), .B2(n3283), .C1(ymem_data1[151]), 
        .C2(n782), .A(n2028), .ZN(n2026) );
  AOI221_X2 U1424 ( .B1(n3234), .B2(ymem_data2[215]), .C1(n3232), .C2(
        ymem_data1[23]), .A(n2031), .ZN(n2030) );
  AOI221_X2 U1426 ( .B1(n3225), .B2(ymem_data1[215]), .C1(n3237), .C2(
        U72_DATA1_23), .A(n2032), .ZN(n2029) );
  OAI22_X2 U1427 ( .A1(n283), .A2(n3198), .B1(n347), .B2(n1815), .ZN(n2032) );
  AOI221_X2 U1430 ( .B1(ymem_data1[214]), .B2(n3283), .C1(ymem_data1[150]), 
        .C2(n782), .A(n2035), .ZN(n2033) );
  AOI221_X2 U1432 ( .B1(n3234), .B2(ymem_data2[214]), .C1(n3232), .C2(
        ymem_data1[22]), .A(n2038), .ZN(n2037) );
  AOI221_X2 U1434 ( .B1(n3225), .B2(ymem_data1[214]), .C1(n3237), .C2(
        U72_DATA1_22), .A(n2039), .ZN(n2036) );
  OAI22_X2 U1435 ( .A1(n284), .A2(n3198), .B1(n348), .B2(n3223), .ZN(n2039) );
  AOI221_X2 U1438 ( .B1(ymem_data1[213]), .B2(n3283), .C1(ymem_data1[149]), 
        .C2(n782), .A(n2042), .ZN(n2040) );
  AOI221_X2 U1440 ( .B1(n3234), .B2(ymem_data2[213]), .C1(n3232), .C2(
        ymem_data1[21]), .A(n2045), .ZN(n2044) );
  AOI221_X2 U1442 ( .B1(n3225), .B2(ymem_data1[213]), .C1(n3237), .C2(
        U72_DATA1_21), .A(n2046), .ZN(n2043) );
  OAI22_X2 U1443 ( .A1(n285), .A2(n3198), .B1(n349), .B2(n1815), .ZN(n2046) );
  AOI221_X2 U1446 ( .B1(ymem_data1[212]), .B2(n3283), .C1(ymem_data1[148]), 
        .C2(n782), .A(n2049), .ZN(n2047) );
  AOI221_X2 U1448 ( .B1(n3234), .B2(ymem_data2[212]), .C1(n3232), .C2(
        ymem_data1[20]), .A(n2052), .ZN(n2051) );
  AOI221_X2 U1450 ( .B1(n3225), .B2(ymem_data1[212]), .C1(n3237), .C2(
        U72_DATA1_20), .A(n2053), .ZN(n2050) );
  OAI22_X2 U1451 ( .A1(n286), .A2(n3198), .B1(n350), .B2(n1815), .ZN(n2053) );
  AOI221_X2 U1456 ( .B1(n3235), .B2(ymem_data2[194]), .C1(n1807), .C2(
        ymem_data1[2]), .A(n2059), .ZN(n2058) );
  AOI221_X2 U1458 ( .B1(n3224), .B2(ymem_data1[194]), .C1(n3237), .C2(
        U72_DATA1_2), .A(n2060), .ZN(n2057) );
  OAI22_X2 U1459 ( .A1(n304), .A2(n3198), .B1(n368), .B2(n1815), .ZN(n2060) );
  AOI221_X2 U1462 ( .B1(ymem_data1[211]), .B2(n3283), .C1(ymem_data1[147]), 
        .C2(n782), .A(n2063), .ZN(n2061) );
  AOI221_X2 U1464 ( .B1(n3235), .B2(ymem_data2[211]), .C1(n1807), .C2(
        ymem_data1[19]), .A(n2066), .ZN(n2065) );
  AOI221_X2 U1466 ( .B1(n3224), .B2(ymem_data1[211]), .C1(n3237), .C2(
        U72_DATA1_19), .A(n2067), .ZN(n2064) );
  OAI22_X2 U1467 ( .A1(n287), .A2(n3198), .B1(n351), .B2(n3223), .ZN(n2067) );
  AOI221_X2 U1470 ( .B1(ymem_data1[210]), .B2(n3283), .C1(ymem_data1[146]), 
        .C2(n782), .A(n2070), .ZN(n2068) );
  AOI221_X2 U1472 ( .B1(n3234), .B2(ymem_data2[210]), .C1(n3232), .C2(
        ymem_data1[18]), .A(n2073), .ZN(n2072) );
  AOI221_X2 U1474 ( .B1(n3224), .B2(ymem_data1[210]), .C1(n3237), .C2(
        U72_DATA1_18), .A(n2074), .ZN(n2071) );
  OAI22_X2 U1475 ( .A1(n288), .A2(n3198), .B1(n352), .B2(n3223), .ZN(n2074) );
  AOI221_X2 U1478 ( .B1(ymem_data1[209]), .B2(n3283), .C1(ymem_data1[145]), 
        .C2(n782), .A(n2077), .ZN(n2075) );
  AOI221_X2 U1480 ( .B1(n3234), .B2(ymem_data2[209]), .C1(n1807), .C2(
        ymem_data1[17]), .A(n2080), .ZN(n2079) );
  AOI221_X2 U1482 ( .B1(n3224), .B2(ymem_data1[209]), .C1(n3237), .C2(
        U72_DATA1_17), .A(n2081), .ZN(n2078) );
  OAI22_X2 U1483 ( .A1(n289), .A2(n3198), .B1(n353), .B2(n3223), .ZN(n2081) );
  AOI221_X2 U1486 ( .B1(ymem_data1[208]), .B2(n3283), .C1(ymem_data1[144]), 
        .C2(n782), .A(n2084), .ZN(n2082) );
  AOI221_X2 U1488 ( .B1(n3234), .B2(ymem_data2[208]), .C1(n3232), .C2(
        ymem_data1[16]), .A(n2087), .ZN(n2086) );
  AOI221_X2 U1490 ( .B1(n3224), .B2(ymem_data1[208]), .C1(n3237), .C2(
        U72_DATA1_16), .A(n2088), .ZN(n2085) );
  OAI22_X2 U1491 ( .A1(n290), .A2(n3198), .B1(n354), .B2(n1815), .ZN(n2088) );
  AOI221_X2 U1496 ( .B1(n3235), .B2(ymem_data2[207]), .C1(n3232), .C2(
        ymem_data1[15]), .A(n2094), .ZN(n2093) );
  AOI221_X2 U1498 ( .B1(n3224), .B2(ymem_data1[207]), .C1(n3237), .C2(
        U72_DATA1_15), .A(n2095), .ZN(n2092) );
  AOI221_X2 U1504 ( .B1(n3234), .B2(ymem_data2[206]), .C1(n3232), .C2(
        ymem_data1[14]), .A(n2101), .ZN(n2100) );
  AOI221_X2 U1506 ( .B1(n3224), .B2(ymem_data1[206]), .C1(n3237), .C2(
        U72_DATA1_14), .A(n2102), .ZN(n2099) );
  OAI22_X2 U1507 ( .A1(n292), .A2(n3198), .B1(n356), .B2(n1815), .ZN(n2102) );
  AOI221_X2 U1510 ( .B1(ymem_data1[205]), .B2(n3283), .C1(ymem_data1[141]), 
        .C2(n782), .A(n2105), .ZN(n2103) );
  AOI221_X2 U1512 ( .B1(n3235), .B2(ymem_data2[205]), .C1(n1807), .C2(
        ymem_data1[13]), .A(n2108), .ZN(n2107) );
  AOI221_X2 U1514 ( .B1(n3224), .B2(ymem_data1[205]), .C1(n3237), .C2(
        U72_DATA1_13), .A(n2109), .ZN(n2106) );
  OAI22_X2 U1515 ( .A1(n293), .A2(n3198), .B1(n357), .B2(n1815), .ZN(n2109) );
  AOI221_X2 U1518 ( .B1(ymem_data1[204]), .B2(n3283), .C1(ymem_data1[140]), 
        .C2(n3280), .A(n2112), .ZN(n2110) );
  AOI221_X2 U1522 ( .B1(n3224), .B2(ymem_data1[204]), .C1(n3236), .C2(
        U72_DATA1_12), .A(n2116), .ZN(n2113) );
  AOI221_X2 U1526 ( .B1(ymem_data1[203]), .B2(n3283), .C1(ymem_data1[139]), 
        .C2(n3280), .A(n2119), .ZN(n2117) );
  AOI221_X2 U1530 ( .B1(n3224), .B2(ymem_data1[203]), .C1(n3236), .C2(
        U72_DATA1_11), .A(n2123), .ZN(n2120) );
  AOI221_X2 U1534 ( .B1(ymem_data1[202]), .B2(n3283), .C1(ymem_data1[138]), 
        .C2(n3280), .A(n2126), .ZN(n2124) );
  AOI221_X2 U1538 ( .B1(n3224), .B2(ymem_data1[202]), .C1(n3237), .C2(
        U72_DATA1_10), .A(n2130), .ZN(n2127) );
  AOI221_X2 U1542 ( .B1(ymem_data1[193]), .B2(n3283), .C1(ymem_data1[129]), 
        .C2(n3280), .A(n2133), .ZN(n2131) );
  AOI221_X2 U1546 ( .B1(n3224), .B2(ymem_data1[193]), .C1(n3236), .C2(
        U72_DATA1_1), .A(n2137), .ZN(n2134) );
  NAND2_X2 U1552 ( .A1(n2140), .A2(n797), .ZN(n628) );
  AOI221_X2 U1553 ( .B1(ymem_data1[192]), .B2(n3283), .C1(ymem_data1[128]), 
        .C2(n3280), .A(n2141), .ZN(n2138) );
  AOI221_X2 U1555 ( .B1(n3235), .B2(ymem_data2[192]), .C1(n1807), .C2(
        ymem_data1[0]), .A(n2144), .ZN(n2143) );
  NAND2_X2 U1557 ( .A1(n813), .A2(exModDone), .ZN(n1811) );
  NAND2_X2 U1559 ( .A1(n1776), .A2(n698), .ZN(n710) );
  NOR2_X2 U1560 ( .A1(n2146), .A2(n107), .ZN(n1776) );
  NAND2_X2 U1561 ( .A1(n780), .A2(exModDone), .ZN(n1810) );
  NOR2_X2 U1562 ( .A1(n852), .A2(n722), .ZN(n780) );
  NAND3_X2 U1563 ( .A1(n690), .A2(n3259), .A3(n737), .ZN(n852) );
  NOR2_X2 U1564 ( .A1(n735), .A2(n132), .ZN(n737) );
  NOR2_X2 U1566 ( .A1(n851), .A2(n722), .ZN(n804) );
  NAND4_X2 U1567 ( .A1(n118), .A2(n88), .A3(n1766), .A4(n3259), .ZN(n851) );
  NOR2_X2 U1568 ( .A1(n1789), .A2(n156), .ZN(n1807) );
  NAND2_X2 U1569 ( .A1(n3262), .A2(n9), .ZN(n1789) );
  NAND2_X2 U1572 ( .A1(n3268), .A2(n9), .ZN(n823) );
  NOR2_X2 U1573 ( .A1(n711), .A2(n2145), .ZN(n849) );
  NAND3_X2 U1574 ( .A1(n1766), .A2(n3259), .A3(n2147), .ZN(n2145) );
  NAND2_X2 U1575 ( .A1(n107), .A2(n698), .ZN(n711) );
  AOI221_X2 U1576 ( .B1(n3224), .B2(ymem_data1[192]), .C1(n3236), .C2(
        U72_DATA1_0), .A(n2148), .ZN(n2142) );
  NAND2_X2 U1578 ( .A1(n805), .A2(exModDone), .ZN(n1815) );
  NOR3_X2 U1579 ( .A1(n95), .A2(n3258), .A3(n1766), .ZN(n854) );
  NOR2_X2 U1581 ( .A1(n857), .A2(n722), .ZN(n812) );
  NAND2_X2 U1582 ( .A1(n95), .A2(n3259), .ZN(n857) );
  NOR2_X2 U1584 ( .A1(n722), .A2(n3259), .ZN(n727) );
  NAND2_X2 U1585 ( .A1(n1791), .A2(n2150), .ZN(U92_Z_0) );
  NOR3_X2 U1587 ( .A1(n829), .A2(exModDone), .A3(yMemDataReadyNextCycle), .ZN(
        n2151) );
  NOR2_X2 U1588 ( .A1(n3204), .A2(n1794), .ZN(n1791) );
  NOR4_X2 U1589 ( .A1(n2152), .A2(n152), .A3(n3300), .A4(exModDone), .ZN(n1794) );
  OAI221_X2 U1590 ( .B1(n179), .B2(n829), .C1(n163), .C2(n3221), .A(n2154), 
        .ZN(U91_Z_9) );
  OAI221_X2 U1591 ( .B1(n180), .B2(n829), .C1(n164), .C2(n3221), .A(n2154), 
        .ZN(U91_Z_8) );
  OAI221_X2 U1592 ( .B1(n181), .B2(n829), .C1(n165), .C2(n3221), .A(n2154), 
        .ZN(U91_Z_7) );
  OAI221_X2 U1593 ( .B1(n182), .B2(n829), .C1(n166), .C2(n3221), .A(n2154), 
        .ZN(U91_Z_6) );
  OAI221_X2 U1594 ( .B1(n183), .B2(n829), .C1(n167), .C2(n3221), .A(n2154), 
        .ZN(U91_Z_5) );
  OAI221_X2 U1595 ( .B1(n184), .B2(n829), .C1(n168), .C2(n3221), .A(n2154), 
        .ZN(U91_Z_4) );
  OAI221_X2 U1596 ( .B1(n185), .B2(n829), .C1(n169), .C2(n3221), .A(n2154), 
        .ZN(U91_Z_3) );
  OAI221_X2 U1597 ( .B1(n186), .B2(n829), .C1(n170), .C2(n3221), .A(n2154), 
        .ZN(U91_Z_2) );
  OAI221_X2 U1598 ( .B1(n173), .B2(n829), .C1(n157), .C2(n3221), .A(n2154), 
        .ZN(U91_Z_15) );
  OAI221_X2 U1599 ( .B1(n174), .B2(n829), .C1(n158), .C2(n3221), .A(n2154), 
        .ZN(U91_Z_14) );
  OAI221_X2 U1600 ( .B1(n175), .B2(n829), .C1(n159), .C2(n3221), .A(n2154), 
        .ZN(U91_Z_13) );
  OAI221_X2 U1601 ( .B1(n176), .B2(n829), .C1(n160), .C2(n3221), .A(n2154), 
        .ZN(U91_Z_12) );
  OAI221_X2 U1602 ( .B1(n177), .B2(n829), .C1(n161), .C2(n3221), .A(n2154), 
        .ZN(U91_Z_11) );
  OAI221_X2 U1603 ( .B1(n178), .B2(n829), .C1(n162), .C2(n3221), .A(n2154), 
        .ZN(U91_Z_10) );
  OAI221_X2 U1604 ( .B1(n187), .B2(n829), .C1(n171), .C2(n3221), .A(n2154), 
        .ZN(U91_Z_1) );
  OAI221_X2 U1605 ( .B1(n188), .B2(n829), .C1(n172), .C2(n3221), .A(n2154), 
        .ZN(U91_Z_0) );
  OAI22_X2 U1608 ( .A1(n133), .A2(n152), .B1(n[2370]), .B2(n1798), .ZN(n831)
         );
  NAND2_X2 U1609 ( .A1(yMemDataReadyNextCycle), .A2(n156), .ZN(n1799) );
  NAND2_X2 U1610 ( .A1(n3219), .A2(n2156), .ZN(n2153) );
  NOR4_X2 U1612 ( .A1(n2159), .A2(n1800), .A3(n3215), .A4(n59), .ZN(n2158) );
  NOR2_X2 U1615 ( .A1(n[2372]), .A2(n[2371]), .ZN(n1798) );
  NOR3_X2 U1616 ( .A1(n722), .A2(n3258), .A3(n688), .ZN(n1800) );
  NAND2_X2 U1617 ( .A1(n2160), .A2(n2161), .ZN(n722) );
  NOR4_X2 U1618 ( .A1(n2162), .A2(n2163), .A3(n2164), .A4(n2165), .ZN(n2161)
         );
  NAND4_X2 U1619 ( .A1(n27), .A2(n26), .A3(n28), .A4(n2166), .ZN(n2165) );
  NOR3_X2 U1620 ( .A1(U72_DATA1_33), .A2(U72_DATA1_35), .A3(U72_DATA1_34), 
        .ZN(n2166) );
  NAND4_X2 U1621 ( .A1(n21), .A2(n20), .A3(n22), .A4(n2167), .ZN(n2164) );
  NOR3_X2 U1622 ( .A1(U72_DATA1_39), .A2(U72_DATA1_40), .A3(U72_DATA1_4), .ZN(
        n2167) );
  NAND4_X2 U1623 ( .A1(n16), .A2(n15), .A3(n17), .A4(n2168), .ZN(n2163) );
  NOR3_X2 U1624 ( .A1(U72_DATA1_44), .A2(U72_DATA1_46), .A3(U72_DATA1_45), 
        .ZN(n2168) );
  NAND4_X2 U1625 ( .A1(n53), .A2(n52), .A3(n11), .A4(n2169), .ZN(n2162) );
  NOR3_X2 U1626 ( .A1(U72_DATA1_7), .A2(U72_DATA1_9), .A3(U72_DATA1_8), .ZN(
        n2169) );
  NOR4_X2 U1627 ( .A1(n2170), .A2(n2171), .A3(n2172), .A4(n2173), .ZN(n2160)
         );
  NAND4_X2 U1628 ( .A1(n57), .A2(n48), .A3(n58), .A4(n2174), .ZN(n2173) );
  NOR3_X2 U1629 ( .A1(U72_DATA1_11), .A2(U72_DATA1_13), .A3(U72_DATA1_12), 
        .ZN(n2174) );
  NAND4_X2 U1630 ( .A1(n43), .A2(n42), .A3(n44), .A4(n2175), .ZN(n2172) );
  NOR3_X2 U1631 ( .A1(U72_DATA1_17), .A2(U72_DATA1_19), .A3(U72_DATA1_18), 
        .ZN(n2175) );
  NAND4_X2 U1632 ( .A1(n38), .A2(n37), .A3(n56), .A4(n2176), .ZN(n2171) );
  NOR3_X2 U1633 ( .A1(U72_DATA1_22), .A2(U72_DATA1_24), .A3(U72_DATA1_23), 
        .ZN(n2176) );
  NAND4_X2 U1634 ( .A1(n32), .A2(n31), .A3(n33), .A4(n2177), .ZN(n2170) );
  NOR3_X2 U1635 ( .A1(U72_DATA1_28), .A2(U72_DATA1_3), .A3(U72_DATA1_29), .ZN(
        n2177) );
  OAI22_X2 U1636 ( .A1(n2178), .A2(n2140), .B1(n3216), .B2(n688), .ZN(n2159)
         );
  NAND2_X2 U1637 ( .A1(n86), .A2(n1771), .ZN(n688) );
  AOI221_X2 U1639 ( .B1(n135), .B2(n690), .C1(n141), .C2(n86), .A(n2179), .ZN(
        n2157) );
  NAND2_X2 U1641 ( .A1(n89), .A2(n728), .ZN(n729) );
  NOR2_X2 U1642 ( .A1(n132), .A2(n111), .ZN(n728) );
  NAND3_X2 U1643 ( .A1(n1771), .A2(n2147), .A3(n1778), .ZN(n2178) );
  NAND2_X2 U1644 ( .A1(n87), .A2(n1766), .ZN(n687) );
  NAND4_X2 U1645 ( .A1(n2182), .A2(n2183), .A3(n2184), .A4(n2185), .ZN(n1766)
         );
  NOR4_X2 U1646 ( .A1(n2186), .A2(n2187), .A3(n2188), .A4(n2189), .ZN(n2185)
         );
  XOR2_X2 U1647 ( .A(n2190), .B(n2191), .Z(n2189) );
  OAI22_X2 U1648 ( .A1(n794), .A2(n447), .B1(n2192), .B2(n319), .ZN(n2191) );
  XOR2_X2 U1649 ( .A(n2193), .B(n2194), .Z(n2188) );
  OAI22_X2 U1650 ( .A1(n794), .A2(n448), .B1(n2192), .B2(n320), .ZN(n2194) );
  XOR2_X2 U1651 ( .A(n2195), .B(n2196), .Z(n2187) );
  OAI22_X2 U1652 ( .A1(n794), .A2(n449), .B1(n2192), .B2(n321), .ZN(n2196) );
  XOR2_X2 U1653 ( .A(n2197), .B(n2198), .Z(n2186) );
  NOR4_X2 U1655 ( .A1(n2199), .A2(n2200), .A3(n2201), .A4(n2202), .ZN(n2184)
         );
  XOR2_X2 U1656 ( .A(n2203), .B(n2204), .Z(n2202) );
  OAI22_X2 U1657 ( .A1(n794), .A2(n443), .B1(n2192), .B2(n315), .ZN(n2204) );
  XOR2_X2 U1658 ( .A(n2205), .B(n2206), .Z(n2201) );
  OAI22_X2 U1659 ( .A1(n794), .A2(n444), .B1(n2192), .B2(n316), .ZN(n2206) );
  XOR2_X2 U1660 ( .A(n2207), .B(n2208), .Z(n2200) );
  OAI22_X2 U1661 ( .A1(n794), .A2(n445), .B1(n2192), .B2(n317), .ZN(n2208) );
  XOR2_X2 U1662 ( .A(n2209), .B(n2210), .Z(n2199) );
  NOR4_X2 U1664 ( .A1(n2211), .A2(n2212), .A3(n2213), .A4(n2214), .ZN(n2183)
         );
  XOR2_X2 U1665 ( .A(n2215), .B(n2216), .Z(n2214) );
  OAI22_X2 U1666 ( .A1(n794), .A2(n439), .B1(n2192), .B2(n311), .ZN(n2216) );
  XOR2_X2 U1667 ( .A(n2217), .B(n2218), .Z(n2213) );
  OAI22_X2 U1668 ( .A1(n794), .A2(n440), .B1(n2192), .B2(n312), .ZN(n2218) );
  XOR2_X2 U1669 ( .A(n2219), .B(n2220), .Z(n2212) );
  OAI22_X2 U1670 ( .A1(n794), .A2(n441), .B1(n2192), .B2(n313), .ZN(n2220) );
  XOR2_X2 U1671 ( .A(n2221), .B(n2222), .Z(n2211) );
  NOR4_X2 U1673 ( .A1(n2223), .A2(n2224), .A3(n2225), .A4(n2226), .ZN(n2182)
         );
  XOR2_X2 U1674 ( .A(n2227), .B(n2228), .Z(n2226) );
  OAI22_X2 U1675 ( .A1(n794), .A2(n435), .B1(n2192), .B2(n307), .ZN(n2228) );
  XOR2_X2 U1676 ( .A(n2229), .B(n2230), .Z(n2225) );
  OAI22_X2 U1677 ( .A1(n794), .A2(n436), .B1(n2192), .B2(n308), .ZN(n2230) );
  XOR2_X2 U1678 ( .A(n2231), .B(n2232), .Z(n2224) );
  XOR2_X2 U1680 ( .A(n2233), .B(n2234), .Z(n2223) );
  OAI22_X2 U1681 ( .A1(n3278), .A2(n438), .B1(n2192), .B2(n310), .ZN(n2234) );
  NAND2_X2 U1683 ( .A1(n88), .A2(n735), .ZN(n2180) );
  NAND4_X2 U1684 ( .A1(n2236), .A2(n2237), .A3(n2238), .A4(n2239), .ZN(n735)
         );
  NOR4_X2 U1685 ( .A1(n2240), .A2(n2241), .A3(n2242), .A4(n2243), .ZN(n2239)
         );
  XNOR2_X2 U1686 ( .A(n2244), .B(n2245), .ZN(n2243) );
  OAI22_X2 U1689 ( .A1(n2235), .A2(n185), .B1(n2248), .B2(n169), .ZN(n2190) );
  XNOR2_X2 U1690 ( .A(n2249), .B(n2250), .ZN(n2242) );
  OAI22_X2 U1693 ( .A1(n2235), .A2(n186), .B1(n2248), .B2(n170), .ZN(n2193) );
  XNOR2_X2 U1694 ( .A(n2251), .B(n2252), .ZN(n2241) );
  OAI22_X2 U1697 ( .A1(n2235), .A2(n187), .B1(n2248), .B2(n171), .ZN(n2195) );
  XNOR2_X2 U1698 ( .A(n2253), .B(n2254), .ZN(n2240) );
  OAI22_X2 U1701 ( .A1(n2235), .A2(n188), .B1(n2248), .B2(n172), .ZN(n2197) );
  NOR4_X2 U1702 ( .A1(n2255), .A2(n2256), .A3(n2257), .A4(n2258), .ZN(n2238)
         );
  XNOR2_X2 U1703 ( .A(n2259), .B(n2260), .ZN(n2258) );
  OAI22_X2 U1706 ( .A1(n2235), .A2(n181), .B1(n2248), .B2(n165), .ZN(n2203) );
  XNOR2_X2 U1707 ( .A(n2261), .B(n2262), .ZN(n2257) );
  OAI22_X2 U1710 ( .A1(n2235), .A2(n182), .B1(n2248), .B2(n166), .ZN(n2205) );
  XNOR2_X2 U1711 ( .A(n2263), .B(n2264), .ZN(n2256) );
  OAI22_X2 U1714 ( .A1(n2235), .A2(n183), .B1(n2248), .B2(n167), .ZN(n2207) );
  XNOR2_X2 U1715 ( .A(n2265), .B(n2266), .ZN(n2255) );
  OAI22_X2 U1718 ( .A1(n2235), .A2(n184), .B1(n2248), .B2(n168), .ZN(n2209) );
  NOR4_X2 U1719 ( .A1(n2267), .A2(n2268), .A3(n2269), .A4(n2270), .ZN(n2237)
         );
  XNOR2_X2 U1720 ( .A(n2271), .B(n2272), .ZN(n2270) );
  OAI22_X2 U1723 ( .A1(n2235), .A2(n177), .B1(n2248), .B2(n161), .ZN(n2215) );
  XNOR2_X2 U1724 ( .A(n2273), .B(n2274), .ZN(n2269) );
  OAI22_X2 U1727 ( .A1(n2235), .A2(n178), .B1(n2248), .B2(n162), .ZN(n2217) );
  XNOR2_X2 U1728 ( .A(n2275), .B(n2276), .ZN(n2268) );
  OAI22_X2 U1731 ( .A1(n2235), .A2(n179), .B1(n2248), .B2(n163), .ZN(n2219) );
  XNOR2_X2 U1732 ( .A(n2277), .B(n2278), .ZN(n2267) );
  OAI22_X2 U1735 ( .A1(n2235), .A2(n180), .B1(n2248), .B2(n164), .ZN(n2221) );
  NOR4_X2 U1736 ( .A1(n2279), .A2(n2280), .A3(n2281), .A4(n2282), .ZN(n2236)
         );
  XNOR2_X2 U1737 ( .A(n2283), .B(n2284), .ZN(n2282) );
  OAI22_X2 U1740 ( .A1(n2235), .A2(n173), .B1(n2248), .B2(n157), .ZN(n2227) );
  XNOR2_X2 U1741 ( .A(n2285), .B(n2286), .ZN(n2281) );
  OAI22_X2 U1744 ( .A1(n2235), .A2(n174), .B1(n2248), .B2(n158), .ZN(n2229) );
  XNOR2_X2 U1745 ( .A(n2287), .B(n2288), .ZN(n2280) );
  OAI22_X2 U1748 ( .A1(n2235), .A2(n175), .B1(n2248), .B2(n159), .ZN(n2231) );
  XNOR2_X2 U1749 ( .A(n2289), .B(n2290), .ZN(n2279) );
  NAND2_X2 U1753 ( .A1(n795), .A2(n791), .ZN(n782) );
  OAI22_X2 U1755 ( .A1(n2235), .A2(n176), .B1(n2248), .B2(n160), .ZN(n2233) );
  NOR2_X2 U1756 ( .A1(n2181), .A2(n118), .ZN(n690) );
  NAND4_X2 U1757 ( .A1(n2292), .A2(n2293), .A3(n2294), .A4(n2295), .ZN(n1771)
         );
  NOR4_X2 U1758 ( .A1(n2296), .A2(n2297), .A3(n2298), .A4(n2299), .ZN(n2295)
         );
  XOR2_X2 U1759 ( .A(n511), .B(n2300), .Z(n2299) );
  XOR2_X2 U1761 ( .A(n512), .B(n2303), .Z(n2298) );
  XOR2_X2 U1763 ( .A(n513), .B(n2304), .Z(n2297) );
  XOR2_X2 U1765 ( .A(n514), .B(n2305), .Z(n2296) );
  NOR4_X2 U1767 ( .A1(n2306), .A2(n2307), .A3(n2308), .A4(n2309), .ZN(n2294)
         );
  XOR2_X2 U1768 ( .A(n507), .B(n2310), .Z(n2309) );
  XOR2_X2 U1770 ( .A(n508), .B(n2311), .Z(n2308) );
  XOR2_X2 U1772 ( .A(n509), .B(n2312), .Z(n2307) );
  XOR2_X2 U1774 ( .A(n510), .B(n2313), .Z(n2306) );
  NOR4_X2 U1776 ( .A1(n2314), .A2(n2315), .A3(n2316), .A4(n2317), .ZN(n2293)
         );
  XOR2_X2 U1777 ( .A(n503), .B(n2318), .Z(n2317) );
  XOR2_X2 U1779 ( .A(n504), .B(n2319), .Z(n2316) );
  XOR2_X2 U1781 ( .A(n505), .B(n2320), .Z(n2315) );
  XOR2_X2 U1783 ( .A(n506), .B(n2321), .Z(n2314) );
  NOR4_X2 U1785 ( .A1(n2322), .A2(n2323), .A3(n2324), .A4(n2325), .ZN(n2292)
         );
  XOR2_X2 U1786 ( .A(n499), .B(n2326), .Z(n2325) );
  XOR2_X2 U1788 ( .A(n500), .B(n2327), .Z(n2324) );
  XOR2_X2 U1790 ( .A(n501), .B(n2328), .Z(n2323) );
  XOR2_X2 U1792 ( .A(n502), .B(n2329), .Z(n2322) );
  NAND3_X2 U1796 ( .A1(n2147), .A2(n698), .A3(n1778), .ZN(n2181) );
  NAND4_X2 U1797 ( .A1(n2330), .A2(n2331), .A3(n2332), .A4(n2333), .ZN(n825)
         );
  NOR4_X2 U1798 ( .A1(n2334), .A2(n2335), .A3(n2336), .A4(n2337), .ZN(n2333)
         );
  XOR2_X2 U1799 ( .A(n2338), .B(n2339), .Z(n2337) );
  OAI22_X2 U1800 ( .A1(n319), .A2(n3278), .B1(n2340), .B2(n447), .ZN(n2339) );
  XOR2_X2 U1801 ( .A(n2341), .B(n2342), .Z(n2336) );
  OAI22_X2 U1802 ( .A1(n320), .A2(n794), .B1(n2340), .B2(n448), .ZN(n2342) );
  XOR2_X2 U1803 ( .A(n2343), .B(n2344), .Z(n2335) );
  OAI22_X2 U1804 ( .A1(n321), .A2(n794), .B1(n2340), .B2(n449), .ZN(n2344) );
  XOR2_X2 U1805 ( .A(n2345), .B(n2346), .Z(n2334) );
  OAI22_X2 U1806 ( .A1(n322), .A2(n794), .B1(n2340), .B2(n450), .ZN(n2346) );
  NOR4_X2 U1807 ( .A1(n2347), .A2(n2348), .A3(n2349), .A4(n2350), .ZN(n2332)
         );
  XOR2_X2 U1808 ( .A(n2351), .B(n2352), .Z(n2350) );
  OAI22_X2 U1809 ( .A1(n315), .A2(n3278), .B1(n2340), .B2(n443), .ZN(n2352) );
  XOR2_X2 U1810 ( .A(n2353), .B(n2354), .Z(n2349) );
  OAI22_X2 U1811 ( .A1(n316), .A2(n794), .B1(n2340), .B2(n444), .ZN(n2354) );
  XOR2_X2 U1812 ( .A(n2355), .B(n2356), .Z(n2348) );
  OAI22_X2 U1813 ( .A1(n317), .A2(n794), .B1(n2340), .B2(n445), .ZN(n2356) );
  XOR2_X2 U1814 ( .A(n2357), .B(n2358), .Z(n2347) );
  OAI22_X2 U1815 ( .A1(n318), .A2(n794), .B1(n2340), .B2(n446), .ZN(n2358) );
  NOR4_X2 U1816 ( .A1(n2359), .A2(n2360), .A3(n2361), .A4(n2362), .ZN(n2331)
         );
  XOR2_X2 U1817 ( .A(n2363), .B(n2364), .Z(n2362) );
  OAI22_X2 U1818 ( .A1(n3278), .A2(n311), .B1(n2340), .B2(n439), .ZN(n2364) );
  XOR2_X2 U1819 ( .A(n2365), .B(n2366), .Z(n2361) );
  OAI22_X2 U1820 ( .A1(n3278), .A2(n312), .B1(n2340), .B2(n440), .ZN(n2366) );
  XOR2_X2 U1821 ( .A(n2367), .B(n2368), .Z(n2360) );
  OAI22_X2 U1822 ( .A1(n3278), .A2(n313), .B1(n2340), .B2(n441), .ZN(n2368) );
  XOR2_X2 U1823 ( .A(n2369), .B(n2373), .Z(n2359) );
  OAI22_X2 U1824 ( .A1(n3278), .A2(n314), .B1(n2340), .B2(n442), .ZN(n2373) );
  NOR4_X2 U1825 ( .A1(n2374), .A2(n2375), .A3(n2376), .A4(n2377), .ZN(n2330)
         );
  XOR2_X2 U1826 ( .A(n2378), .B(n2379), .Z(n2377) );
  OAI22_X2 U1827 ( .A1(n307), .A2(n794), .B1(n2340), .B2(n435), .ZN(n2379) );
  XOR2_X2 U1828 ( .A(n2380), .B(n2381), .Z(n2376) );
  OAI22_X2 U1829 ( .A1(n308), .A2(n794), .B1(n2340), .B2(n436), .ZN(n2381) );
  XOR2_X2 U1830 ( .A(n2382), .B(n2383), .Z(n2375) );
  OAI22_X2 U1831 ( .A1(n309), .A2(n794), .B1(n2340), .B2(n437), .ZN(n2383) );
  XOR2_X2 U1832 ( .A(n2384), .B(n2385), .Z(n2374) );
  OAI22_X2 U1833 ( .A1(n3278), .A2(n310), .B1(n2340), .B2(n438), .ZN(n2385) );
  NAND4_X2 U1834 ( .A1(n2388), .A2(n2389), .A3(n2390), .A4(n2391), .ZN(n2146)
         );
  NOR4_X2 U1835 ( .A1(n2392), .A2(n2393), .A3(n2394), .A4(n2395), .ZN(n2391)
         );
  XOR2_X2 U1836 ( .A(n2338), .B(ymem_data2[179]), .Z(n2395) );
  XOR2_X2 U1837 ( .A(n2341), .B(ymem_data2[178]), .Z(n2394) );
  XOR2_X2 U1838 ( .A(n2343), .B(ymem_data2[177]), .Z(n2393) );
  XOR2_X2 U1839 ( .A(n2345), .B(ymem_data2[176]), .Z(n2392) );
  NOR4_X2 U1840 ( .A1(n2396), .A2(n2397), .A3(n2398), .A4(n2399), .ZN(n2390)
         );
  XOR2_X2 U1841 ( .A(n2351), .B(ymem_data2[183]), .Z(n2399) );
  XOR2_X2 U1842 ( .A(n2353), .B(ymem_data2[182]), .Z(n2398) );
  XOR2_X2 U1843 ( .A(n2355), .B(ymem_data2[181]), .Z(n2397) );
  XOR2_X2 U1844 ( .A(n2357), .B(ymem_data2[180]), .Z(n2396) );
  NOR4_X2 U1845 ( .A1(n2400), .A2(n2401), .A3(n2402), .A4(n2403), .ZN(n2389)
         );
  XOR2_X2 U1846 ( .A(n2363), .B(ymem_data2[187]), .Z(n2403) );
  XOR2_X2 U1847 ( .A(n2365), .B(ymem_data2[186]), .Z(n2402) );
  XOR2_X2 U1848 ( .A(n2367), .B(ymem_data2[185]), .Z(n2401) );
  XOR2_X2 U1849 ( .A(n2369), .B(ymem_data2[184]), .Z(n2400) );
  NOR4_X2 U1850 ( .A1(n2404), .A2(n2405), .A3(n2406), .A4(n2407), .ZN(n2388)
         );
  XOR2_X2 U1851 ( .A(n2378), .B(ymem_data2[191]), .Z(n2407) );
  XOR2_X2 U1852 ( .A(n2380), .B(ymem_data2[190]), .Z(n2406) );
  XOR2_X2 U1853 ( .A(n2382), .B(ymem_data2[189]), .Z(n2405) );
  XOR2_X2 U1854 ( .A(n2384), .B(ymem_data2[188]), .Z(n2404) );
  NAND4_X2 U1855 ( .A1(n2408), .A2(n2409), .A3(n2410), .A4(n2411), .ZN(n698)
         );
  NOR4_X2 U1856 ( .A1(n2412), .A2(n2413), .A3(n2414), .A4(n2415), .ZN(n2411)
         );
  XOR2_X2 U1857 ( .A(n2416), .B(n2417), .Z(n2415) );
  OAI22_X2 U1858 ( .A1(n2418), .A2(n511), .B1(n2419), .B2(n383), .ZN(n2417) );
  OAI22_X2 U1859 ( .A1(n3205), .A2(n185), .B1(n2420), .B2(n169), .ZN(n2416) );
  XOR2_X2 U1860 ( .A(n2421), .B(n2422), .Z(n2414) );
  OAI22_X2 U1861 ( .A1(n2418), .A2(n512), .B1(n2419), .B2(n384), .ZN(n2422) );
  OAI22_X2 U1862 ( .A1(n3205), .A2(n186), .B1(n2420), .B2(n170), .ZN(n2421) );
  XOR2_X2 U1863 ( .A(n2423), .B(n2424), .Z(n2413) );
  OAI22_X2 U1864 ( .A1(n2418), .A2(n513), .B1(n2419), .B2(n385), .ZN(n2424) );
  OAI22_X2 U1865 ( .A1(n3205), .A2(n187), .B1(n2420), .B2(n171), .ZN(n2423) );
  XOR2_X2 U1866 ( .A(n2425), .B(n2426), .Z(n2412) );
  OAI22_X2 U1867 ( .A1(n2418), .A2(n514), .B1(n2419), .B2(n386), .ZN(n2426) );
  OAI22_X2 U1868 ( .A1(n3205), .A2(n188), .B1(n2420), .B2(n172), .ZN(n2425) );
  NOR4_X2 U1869 ( .A1(n2427), .A2(n2428), .A3(n2429), .A4(n2430), .ZN(n2410)
         );
  XOR2_X2 U1870 ( .A(n2431), .B(n2432), .Z(n2430) );
  OAI22_X2 U1871 ( .A1(n2418), .A2(n507), .B1(n2419), .B2(n379), .ZN(n2432) );
  OAI22_X2 U1872 ( .A1(n3205), .A2(n181), .B1(n2420), .B2(n165), .ZN(n2431) );
  XOR2_X2 U1873 ( .A(n2433), .B(n2434), .Z(n2429) );
  OAI22_X2 U1874 ( .A1(n2418), .A2(n508), .B1(n2419), .B2(n380), .ZN(n2434) );
  OAI22_X2 U1875 ( .A1(n3205), .A2(n182), .B1(n2420), .B2(n166), .ZN(n2433) );
  XOR2_X2 U1876 ( .A(n2435), .B(n2436), .Z(n2428) );
  OAI22_X2 U1877 ( .A1(n2418), .A2(n509), .B1(n2419), .B2(n381), .ZN(n2436) );
  OAI22_X2 U1878 ( .A1(n3205), .A2(n183), .B1(n2420), .B2(n167), .ZN(n2435) );
  XOR2_X2 U1879 ( .A(n2437), .B(n2438), .Z(n2427) );
  OAI22_X2 U1880 ( .A1(n2418), .A2(n510), .B1(n2419), .B2(n382), .ZN(n2438) );
  OAI22_X2 U1881 ( .A1(n3205), .A2(n184), .B1(n2420), .B2(n168), .ZN(n2437) );
  NOR4_X2 U1882 ( .A1(n2439), .A2(n2440), .A3(n2441), .A4(n2442), .ZN(n2409)
         );
  XOR2_X2 U1883 ( .A(n2443), .B(n2444), .Z(n2442) );
  OAI22_X2 U1884 ( .A1(n2418), .A2(n503), .B1(n2419), .B2(n375), .ZN(n2444) );
  OAI22_X2 U1885 ( .A1(n3205), .A2(n177), .B1(n2420), .B2(n161), .ZN(n2443) );
  XOR2_X2 U1886 ( .A(n2445), .B(n2446), .Z(n2441) );
  OAI22_X2 U1887 ( .A1(n2418), .A2(n504), .B1(n2419), .B2(n376), .ZN(n2446) );
  OAI22_X2 U1888 ( .A1(n3205), .A2(n178), .B1(n2420), .B2(n162), .ZN(n2445) );
  XOR2_X2 U1889 ( .A(n2447), .B(n2448), .Z(n2440) );
  OAI22_X2 U1890 ( .A1(n2418), .A2(n505), .B1(n2419), .B2(n377), .ZN(n2448) );
  OAI22_X2 U1891 ( .A1(n3205), .A2(n179), .B1(n2420), .B2(n163), .ZN(n2447) );
  XOR2_X2 U1892 ( .A(n2449), .B(n2450), .Z(n2439) );
  OAI22_X2 U1893 ( .A1(n2418), .A2(n506), .B1(n2419), .B2(n378), .ZN(n2450) );
  OAI22_X2 U1894 ( .A1(n3205), .A2(n180), .B1(n2420), .B2(n164), .ZN(n2449) );
  NOR4_X2 U1895 ( .A1(n2451), .A2(n2452), .A3(n2453), .A4(n2454), .ZN(n2408)
         );
  XOR2_X2 U1896 ( .A(n2455), .B(n2456), .Z(n2454) );
  OAI22_X2 U1897 ( .A1(n2418), .A2(n499), .B1(n2419), .B2(n371), .ZN(n2456) );
  OAI22_X2 U1898 ( .A1(n3205), .A2(n173), .B1(n2420), .B2(n157), .ZN(n2455) );
  XOR2_X2 U1899 ( .A(n2457), .B(n2458), .Z(n2453) );
  OAI22_X2 U1900 ( .A1(n2418), .A2(n500), .B1(n2419), .B2(n372), .ZN(n2458) );
  OAI22_X2 U1901 ( .A1(n3205), .A2(n174), .B1(n2420), .B2(n158), .ZN(n2457) );
  XOR2_X2 U1902 ( .A(n2459), .B(n2460), .Z(n2452) );
  OAI22_X2 U1903 ( .A1(n2418), .A2(n501), .B1(n2419), .B2(n373), .ZN(n2460) );
  OAI22_X2 U1904 ( .A1(n3205), .A2(n175), .B1(n2420), .B2(n159), .ZN(n2459) );
  XOR2_X2 U1905 ( .A(n2461), .B(n2462), .Z(n2451) );
  OAI22_X2 U1906 ( .A1(n2418), .A2(n502), .B1(n2419), .B2(n374), .ZN(n2462) );
  NAND3_X2 U1908 ( .A1(n793), .A2(n776), .A3(n3286), .ZN(n2302) );
  OAI22_X2 U1910 ( .A1(n3205), .A2(n176), .B1(n2420), .B2(n160), .ZN(n2461) );
  NAND2_X2 U1912 ( .A1(n717), .A2(n3278), .ZN(n2291) );
  NAND4_X2 U1913 ( .A1(n2463), .A2(n2464), .A3(n2465), .A4(n2466), .ZN(n2147)
         );
  NOR4_X2 U1914 ( .A1(n2467), .A2(n2468), .A3(n2469), .A4(n2470), .ZN(n2466)
         );
  XNOR2_X2 U1915 ( .A(n2338), .B(n2471), .ZN(n2470) );
  OAI22_X2 U1917 ( .A1(n2473), .A2(n169), .B1(n3205), .B2(n185), .ZN(n2338) );
  XNOR2_X2 U1918 ( .A(n2341), .B(n2474), .ZN(n2469) );
  OAI22_X2 U1920 ( .A1(n2473), .A2(n170), .B1(n3205), .B2(n186), .ZN(n2341) );
  XNOR2_X2 U1921 ( .A(n2343), .B(n2475), .ZN(n2468) );
  OAI22_X2 U1923 ( .A1(n2473), .A2(n171), .B1(n3205), .B2(n187), .ZN(n2343) );
  XNOR2_X2 U1924 ( .A(n2345), .B(n2476), .ZN(n2467) );
  OAI22_X2 U1926 ( .A1(n2473), .A2(n172), .B1(n3205), .B2(n188), .ZN(n2345) );
  NOR4_X2 U1927 ( .A1(n2477), .A2(n2478), .A3(n2479), .A4(n2480), .ZN(n2465)
         );
  XNOR2_X2 U1928 ( .A(n2351), .B(n2481), .ZN(n2480) );
  OAI22_X2 U1930 ( .A1(n2473), .A2(n165), .B1(n3205), .B2(n181), .ZN(n2351) );
  XNOR2_X2 U1931 ( .A(n2353), .B(n2482), .ZN(n2479) );
  OAI22_X2 U1933 ( .A1(n2473), .A2(n166), .B1(n3205), .B2(n182), .ZN(n2353) );
  XNOR2_X2 U1934 ( .A(n2355), .B(n2483), .ZN(n2478) );
  OAI22_X2 U1936 ( .A1(n2473), .A2(n167), .B1(n3205), .B2(n183), .ZN(n2355) );
  XNOR2_X2 U1937 ( .A(n2357), .B(n2484), .ZN(n2477) );
  OAI22_X2 U1939 ( .A1(n2473), .A2(n168), .B1(n3205), .B2(n184), .ZN(n2357) );
  NOR4_X2 U1940 ( .A1(n2485), .A2(n2486), .A3(n2487), .A4(n2488), .ZN(n2464)
         );
  XNOR2_X2 U1941 ( .A(n2363), .B(n2489), .ZN(n2488) );
  OAI22_X2 U1943 ( .A1(n2473), .A2(n161), .B1(n3205), .B2(n177), .ZN(n2363) );
  XNOR2_X2 U1944 ( .A(n2365), .B(n2490), .ZN(n2487) );
  OAI22_X2 U1946 ( .A1(n2473), .A2(n162), .B1(n3205), .B2(n178), .ZN(n2365) );
  XNOR2_X2 U1947 ( .A(n2367), .B(n2491), .ZN(n2486) );
  OAI22_X2 U1949 ( .A1(n2473), .A2(n163), .B1(n3205), .B2(n179), .ZN(n2367) );
  XNOR2_X2 U1950 ( .A(n2369), .B(n2492), .ZN(n2485) );
  OAI22_X2 U1952 ( .A1(n2473), .A2(n164), .B1(n3205), .B2(n180), .ZN(n2369) );
  NOR4_X2 U1953 ( .A1(n2493), .A2(n2494), .A3(n2495), .A4(n2496), .ZN(n2463)
         );
  XNOR2_X2 U1954 ( .A(n2378), .B(n2497), .ZN(n2496) );
  OAI22_X2 U1956 ( .A1(n2473), .A2(n157), .B1(n3205), .B2(n173), .ZN(n2378) );
  XNOR2_X2 U1957 ( .A(n2380), .B(n2498), .ZN(n2495) );
  OAI22_X2 U1959 ( .A1(n2473), .A2(n158), .B1(n3205), .B2(n174), .ZN(n2380) );
  XNOR2_X2 U1960 ( .A(n2382), .B(n2499), .ZN(n2494) );
  OAI22_X2 U1962 ( .A1(n2473), .A2(n159), .B1(n3205), .B2(n175), .ZN(n2382) );
  XNOR2_X2 U1963 ( .A(n2384), .B(n2500), .ZN(n2493) );
  OAI22_X2 U1966 ( .A1(n2473), .A2(n160), .B1(n3205), .B2(n176), .ZN(n2384) );
  NOR2_X2 U1967 ( .A1(n121), .A2(n135), .ZN(n2501) );
  NAND2_X2 U1968 ( .A1(n122), .A2(n3291), .ZN(n797) );
  NAND3_X2 U1969 ( .A1(n138), .A2(n2502), .A3(n693), .ZN(n701) );
  NAND2_X2 U1971 ( .A1(n3220), .A2(n3291), .ZN(n791) );
  NAND2_X2 U1972 ( .A1(n146), .A2(n3291), .ZN(n793) );
  NAND2_X2 U1973 ( .A1(n146), .A2(n150), .ZN(n794) );
  NOR4_X2 U1974 ( .A1(n130), .A2(n113), .A3(n117), .A4(n139), .ZN(n2387) );
  NAND2_X2 U1975 ( .A1(n3220), .A2(n150), .ZN(n795) );
  NAND2_X2 U1977 ( .A1(n120), .A2(n150), .ZN(n2140) );
  NAND3_X2 U1978 ( .A1(n138), .A2(n2505), .A3(n732), .ZN(n739) );
  NOR3_X2 U1979 ( .A1(n372), .A2(n373), .A3(n371), .ZN(n2503) );
  NAND2_X2 U1980 ( .A1(n115), .A2(n150), .ZN(n775) );
  NAND2_X2 U1981 ( .A1(n116), .A2(n138), .ZN(n734) );
  NAND2_X2 U1982 ( .A1(n2507), .A2(n3258), .ZN(n2505) );
  NAND3_X2 U1983 ( .A1(n2508), .A2(n2509), .A3(n2510), .ZN(n856) );
  NOR4_X2 U1984 ( .A1(n2511), .A2(n2512), .A3(n2513), .A4(n2514), .ZN(n2510)
         );
  XOR2_X2 U1985 ( .A(n2515), .B(n2516), .Z(n2514) );
  AOI221_X2 U1987 ( .B1(chng_col[3]), .B2(n3287), .C1(chng_row[3]), .C2(n130), 
        .A(n2517), .ZN(n2515) );
  XOR2_X2 U1988 ( .A(n2518), .B(n2519), .Z(n2513) );
  AOI221_X2 U1990 ( .B1(chng_col[2]), .B2(n3287), .C1(chng_row[2]), .C2(n130), 
        .A(n2520), .ZN(n2518) );
  XOR2_X2 U1992 ( .A(n2523), .B(n2524), .Z(n2522) );
  OAI221_X2 U1994 ( .B1(n3286), .B2(n188), .C1(n717), .C2(n172), .A(n2525), 
        .ZN(n2523) );
  XOR2_X2 U1995 ( .A(n2526), .B(n2527), .Z(n2521) );
  OAI221_X2 U1997 ( .B1(n187), .B2(n3286), .C1(n171), .C2(n717), .A(n2528), 
        .ZN(n2526) );
  NAND4_X2 U1998 ( .A1(n2530), .A2(n2531), .A3(n2532), .A4(n2533), .ZN(n2511)
         );
  XOR2_X2 U1999 ( .A(n2534), .B(n2535), .Z(n2533) );
  OAI221_X2 U2001 ( .B1(n3286), .B2(n184), .C1(n717), .C2(n168), .A(n2536), 
        .ZN(n2534) );
  XOR2_X2 U2002 ( .A(n2537), .B(n2538), .Z(n2532) );
  OAI221_X2 U2004 ( .B1(n3286), .B2(n183), .C1(n717), .C2(n167), .A(n2539), 
        .ZN(n2537) );
  XOR2_X2 U2005 ( .A(n2540), .B(n2541), .Z(n2531) );
  OAI221_X2 U2007 ( .B1(n3286), .B2(n182), .C1(n717), .C2(n166), .A(n2542), 
        .ZN(n2540) );
  XOR2_X2 U2008 ( .A(n2543), .B(n2544), .Z(n2530) );
  OAI221_X2 U2010 ( .B1(n3286), .B2(n181), .C1(n717), .C2(n165), .A(n2545), 
        .ZN(n2543) );
  AOI221_X2 U2011 ( .B1(n2546), .B2(n194), .C1(n2547), .C2(n193), .A(n2548), 
        .ZN(n2509) );
  OAI221_X2 U2012 ( .B1(n131), .B2(n2549), .C1(ymem_data1[248]), .C2(n128), 
        .A(n2550), .ZN(n2548) );
  NOR2_X2 U2014 ( .A1(n2558), .A2(n2559), .ZN(n2549) );
  OAI221_X2 U2015 ( .B1(n2553), .B2(n190), .C1(n2529), .C2(n189), .A(n2560), 
        .ZN(n2559) );
  OAI22_X2 U2017 ( .A1(n2561), .A2(n173), .B1(n2562), .B2(n157), .ZN(n2529) );
  OAI221_X2 U2018 ( .B1(n2547), .B2(n193), .C1(n2556), .C2(n192), .A(n2563), 
        .ZN(n2558) );
  OAI22_X2 U2020 ( .A1(n2561), .A2(n180), .B1(n2562), .B2(n164), .ZN(n2557) );
  OAI22_X2 U2022 ( .A1(n2561), .A2(n178), .B1(n2562), .B2(n162), .ZN(n2547) );
  OAI22_X2 U2023 ( .A1(n2561), .A2(n179), .B1(n2562), .B2(n163), .ZN(n2546) );
  AOI221_X2 U2024 ( .B1(n2554), .B2(n191), .C1(n2553), .C2(n190), .A(n2564), 
        .ZN(n2508) );
  OAI22_X2 U2025 ( .A1(ymem_data1[252]), .A2(n125), .B1(ymem_data1[251]), .B2(
        n126), .ZN(n2564) );
  OAI22_X2 U2026 ( .A1(n2561), .A2(n177), .B1(n2562), .B2(n161), .ZN(n2556) );
  OAI22_X2 U2027 ( .A1(n2561), .A2(n176), .B1(n2562), .B2(n160), .ZN(n2555) );
  OAI22_X2 U2028 ( .A1(n2561), .A2(n174), .B1(n2562), .B2(n158), .ZN(n2553) );
  OAI22_X2 U2029 ( .A1(n2561), .A2(n175), .B1(n2562), .B2(n159), .ZN(n2554) );
  NOR2_X2 U2030 ( .A1(n3291), .A2(n130), .ZN(n2562) );
  NOR2_X2 U2031 ( .A1(n150), .A2(n3287), .ZN(n2561) );
  NAND3_X2 U2032 ( .A1(n[2370]), .A2(n149), .A3(n[2371]), .ZN(n715) );
  NAND2_X2 U2033 ( .A1(n133), .A2(n152), .ZN(n717) );
  NAND2_X2 U2034 ( .A1(n[2371]), .A2(n[2372]), .ZN(n2152) );
  NAND2_X2 U2035 ( .A1(n136), .A2(n3291), .ZN(n776) );
  NAND2_X2 U2036 ( .A1(n137), .A2(n138), .ZN(n697) );
  NAND2_X2 U2037 ( .A1(n2504), .A2(n695), .ZN(n692) );
  NAND4_X2 U2038 ( .A1(n2565), .A2(n2566), .A3(n2567), .A4(n2568), .ZN(n695)
         );
  NOR3_X2 U2039 ( .A1(n2569), .A2(n2570), .A3(n2571), .ZN(n2568) );
  XNOR2_X2 U2040 ( .A(n2525), .B(ymem_data1[240]), .ZN(n2571) );
  XNOR2_X2 U2041 ( .A(n2528), .B(ymem_data1[241]), .ZN(n2570) );
  XNOR2_X2 U2042 ( .A(n2536), .B(ymem_data1[244]), .ZN(n2569) );
  NOR3_X2 U2043 ( .A1(n2572), .A2(n2573), .A3(n2574), .ZN(n2567) );
  XOR2_X2 U2044 ( .A(n2517), .B(ymem_data1[243]), .Z(n2574) );
  XOR2_X2 U2045 ( .A(n2520), .B(ymem_data1[242]), .Z(n2573) );
  XNOR2_X2 U2046 ( .A(n2545), .B(ymem_data1[247]), .ZN(n2572) );
  NOR3_X2 U2047 ( .A1(n191), .A2(n2575), .A3(n2576), .ZN(n2566) );
  XNOR2_X2 U2048 ( .A(n2542), .B(ymem_data1[246]), .ZN(n2576) );
  XNOR2_X2 U2049 ( .A(n2539), .B(ymem_data1[245]), .ZN(n2575) );
  NOR3_X2 U2050 ( .A1(n2577), .A2(n190), .A3(n189), .ZN(n2565) );
  NAND4_X2 U2051 ( .A1(n2578), .A2(n2579), .A3(n2580), .A4(n2581), .ZN(n2504)
         );
  NOR3_X2 U2052 ( .A1(n2582), .A2(n2583), .A3(n2584), .ZN(n2581) );
  XOR2_X2 U2053 ( .A(n2525), .B(n258), .Z(n2584) );
  XOR2_X2 U2054 ( .A(n2528), .B(n257), .Z(n2583) );
  XOR2_X2 U2055 ( .A(n2536), .B(n254), .Z(n2582) );
  NOR3_X2 U2056 ( .A1(n2585), .A2(n2586), .A3(n2587), .ZN(n2580) );
  XOR2_X2 U2057 ( .A(n2517), .B(ymem_data1[179]), .Z(n2587) );
  XOR2_X2 U2058 ( .A(n2520), .B(ymem_data1[178]), .Z(n2586) );
  XOR2_X2 U2059 ( .A(n2545), .B(n251), .Z(n2585) );
  NOR3_X2 U2060 ( .A1(n2577), .A2(n2588), .A3(n2589), .ZN(n2579) );
  XOR2_X2 U2061 ( .A(n2542), .B(n252), .Z(n2589) );
  XOR2_X2 U2062 ( .A(n2539), .B(n253), .Z(n2588) );
  NOR3_X2 U2063 ( .A1(n243), .A2(n245), .A3(n244), .ZN(n2578) );
  NAND2_X2 U2064 ( .A1(n2507), .A2(n2506), .ZN(n2502) );
  AND4_X2 U2065 ( .A1(n2590), .A2(n2591), .A3(n2592), .A4(n2593), .ZN(n2506)
         );
  NOR4_X2 U2066 ( .A1(n2594), .A2(n2595), .A3(n2596), .A4(n2597), .ZN(n2593)
         );
  XNOR2_X2 U2067 ( .A(n2545), .B(n2598), .ZN(n2597) );
  OAI22_X2 U2068 ( .A1(n3218), .A2(n379), .B1(n2156), .B2(n315), .ZN(n2598) );
  XNOR2_X2 U2070 ( .A(n2542), .B(n2599), .ZN(n2596) );
  OAI22_X2 U2071 ( .A1(n634), .A2(n380), .B1(n2156), .B2(n316), .ZN(n2599) );
  XNOR2_X2 U2073 ( .A(n2539), .B(n2600), .ZN(n2595) );
  OAI22_X2 U2074 ( .A1(n634), .A2(n381), .B1(n2156), .B2(n317), .ZN(n2600) );
  XNOR2_X2 U2076 ( .A(n2536), .B(n2601), .ZN(n2594) );
  OAI22_X2 U2077 ( .A1(n634), .A2(n382), .B1(n2156), .B2(n318), .ZN(n2601) );
  NOR3_X2 U2079 ( .A1(n2602), .A2(n2577), .A3(n2603), .ZN(n2592) );
  XNOR2_X2 U2080 ( .A(n2528), .B(n2604), .ZN(n2603) );
  OAI22_X2 U2081 ( .A1(n634), .A2(n385), .B1(n2156), .B2(n321), .ZN(n2604) );
  OAI22_X2 U2083 ( .A1(n2605), .A2(n3218), .B1(n2606), .B2(n2156), .ZN(n2577)
         );
  NOR2_X2 U2084 ( .A1(n2607), .A2(n2608), .ZN(n2606) );
  NAND4_X2 U2085 ( .A1(n162), .A2(n161), .A3(n160), .A4(n159), .ZN(n2608) );
  NAND4_X2 U2086 ( .A1(n158), .A2(n157), .A3(n164), .A4(n163), .ZN(n2607) );
  NOR2_X2 U2087 ( .A1(n2609), .A2(n2610), .ZN(n2605) );
  NAND4_X2 U2088 ( .A1(n178), .A2(n177), .A3(n176), .A4(n175), .ZN(n2610) );
  NAND4_X2 U2089 ( .A1(n174), .A2(n173), .A3(n180), .A4(n179), .ZN(n2609) );
  XNOR2_X2 U2090 ( .A(n2525), .B(n2611), .ZN(n2602) );
  OAI22_X2 U2091 ( .A1(n634), .A2(n386), .B1(n2156), .B2(n322), .ZN(n2611) );
  XOR2_X2 U2093 ( .A(n2520), .B(n2612), .Z(n2591) );
  OAI22_X2 U2095 ( .A1(n3219), .A2(n186), .B1(n2156), .B2(n170), .ZN(n2520) );
  XOR2_X2 U2096 ( .A(n2517), .B(n2613), .Z(n2590) );
  OAI22_X2 U2098 ( .A1(n3219), .A2(n185), .B1(n2156), .B2(n169), .ZN(n2517) );
  NAND3_X2 U2100 ( .A1(n[2370]), .A2(n151), .A3(n[2372]), .ZN(n634) );
  NOR3_X2 U2101 ( .A1(n308), .A2(n309), .A3(n307), .ZN(n2507) );
  INV_X4 U2102 ( .A(n766), .ZN(n1) );
  INV_X4 U2103 ( .A(n1792), .ZN(n2) );
  INV_X4 U2104 ( .A(n1800), .ZN(n3) );
  INV_X4 U2105 ( .A(n823), .ZN(n4) );
  INV_X4 U2106 ( .A(n1789), .ZN(n5) );
  INV_X4 U2107 ( .A(n811), .ZN(n6) );
  INV_X4 U2109 ( .A(n786), .ZN(n8) );
  INV_X4 U2110 ( .A(n722), .ZN(n9) );
  INV_X4 U2111 ( .A(n798), .ZN(n10) );
  INV_X4 U2112 ( .A(n829), .ZN(n59) );
  INV_X4 U2113 ( .A(n763), .ZN(n60) );
  INV_X4 U2114 ( .A(n762), .ZN(n61) );
  INV_X4 U2115 ( .A(n761), .ZN(n62) );
  INV_X4 U2116 ( .A(n760), .ZN(n63) );
  INV_X4 U2117 ( .A(n759), .ZN(n64) );
  INV_X4 U2118 ( .A(n758), .ZN(n65) );
  INV_X4 U2119 ( .A(n757), .ZN(n66) );
  INV_X4 U2120 ( .A(n756), .ZN(n67) );
  INV_X4 U2121 ( .A(n755), .ZN(n68) );
  INV_X4 U2122 ( .A(n754), .ZN(n69) );
  INV_X4 U2123 ( .A(n753), .ZN(n70) );
  INV_X4 U2124 ( .A(n627), .ZN(n71) );
  INV_X4 U2126 ( .A(n629), .ZN(n73) );
  INV_X4 U2128 ( .A(n686), .ZN(n75) );
  INV_X4 U2129 ( .A(n682), .ZN(n76) );
  INV_X4 U2130 ( .A(n678), .ZN(n77) );
  INV_X4 U2131 ( .A(n674), .ZN(n78) );
  INV_X4 U2132 ( .A(n670), .ZN(n79) );
  INV_X4 U2133 ( .A(n666), .ZN(n80) );
  INV_X4 U2134 ( .A(n662), .ZN(n81) );
  INV_X4 U2135 ( .A(n658), .ZN(n82) );
  INV_X4 U2136 ( .A(n654), .ZN(n83) );
  INV_X4 U2137 ( .A(n650), .ZN(n84) );
  INV_X4 U2138 ( .A(n638), .ZN(n85) );
  INV_X4 U2139 ( .A(n687), .ZN(n86) );
  INV_X4 U2140 ( .A(n2180), .ZN(n87) );
  INV_X4 U2141 ( .A(n2181), .ZN(n88) );
  INV_X4 U2142 ( .A(n2178), .ZN(n89) );
  INV_X4 U2143 ( .A(n743), .ZN(n90) );
  INV_X4 U2144 ( .A(n1783), .ZN(n91) );
  INV_X4 U2146 ( .A(n784), .ZN(n93) );
  INV_X4 U2147 ( .A(n1769), .ZN(n94) );
  INV_X4 U2148 ( .A(n2147), .ZN(n95) );
  INV_X4 U2149 ( .A(n751), .ZN(n96) );
  INV_X4 U2150 ( .A(n706), .ZN(n97) );
  INV_X4 U2151 ( .A(n749), .ZN(n98) );
  INV_X4 U2152 ( .A(n1775), .ZN(n99) );
  INV_X4 U2153 ( .A(n814), .ZN(n100) );
  INV_X4 U2154 ( .A(n745), .ZN(n101) );
  INV_X4 U2155 ( .A(n1776), .ZN(n102) );
  INV_X4 U2158 ( .A(n748), .ZN(n105) );
  INV_X4 U2160 ( .A(n825), .ZN(n107) );
  INV_X4 U2162 ( .A(n698), .ZN(n109) );
  INV_X4 U2163 ( .A(n815), .ZN(n110) );
  INV_X4 U2164 ( .A(n735), .ZN(n111) );
  INV_X4 U2165 ( .A(n792), .ZN(n112) );
  INV_X4 U2168 ( .A(n734), .ZN(n115) );
  INV_X4 U2169 ( .A(n2505), .ZN(n116) );
  INV_X4 U2170 ( .A(n2140), .ZN(n117) );
  INV_X4 U2171 ( .A(n1771), .ZN(n118) );
  INV_X4 U2173 ( .A(n739), .ZN(n120) );
  INV_X4 U2174 ( .A(n797), .ZN(n121) );
  INV_X4 U2175 ( .A(n701), .ZN(n122) );
  INV_X4 U2177 ( .A(n2554), .ZN(n124) );
  INV_X4 U2178 ( .A(n2555), .ZN(n125) );
  INV_X4 U2179 ( .A(n2556), .ZN(n126) );
  INV_X4 U2180 ( .A(n2546), .ZN(n127) );
  INV_X4 U2181 ( .A(n2557), .ZN(n128) );
  INV_X4 U2182 ( .A(n2529), .ZN(n129) );
  INV_X4 U2184 ( .A(n765), .ZN(n131) );
  INV_X4 U2186 ( .A(n2152), .ZN(n133) );
  INV_X4 U2187 ( .A(n1794), .ZN(n134) );
  INV_X4 U2188 ( .A(n776), .ZN(n135) );
  INV_X4 U2189 ( .A(n697), .ZN(n136) );
  INV_X4 U2190 ( .A(n2502), .ZN(n137) );
  INV_X4 U2191 ( .A(n692), .ZN(n138) );
  INV_X4 U2192 ( .A(n795), .ZN(n139) );
  INV_X4 U2194 ( .A(n791), .ZN(n141) );
  INV_X4 U2198 ( .A(n793), .ZN(n145) );
  INV_X4 U2204 ( .A(exModDone), .ZN(n156) );
  INV_X4 U2205 ( .A(chng_row[15]), .ZN(n157) );
  INV_X4 U2206 ( .A(chng_row[14]), .ZN(n158) );
  INV_X4 U2207 ( .A(chng_row[13]), .ZN(n159) );
  INV_X4 U2208 ( .A(chng_row[12]), .ZN(n160) );
  INV_X4 U2209 ( .A(chng_row[11]), .ZN(n161) );
  INV_X4 U2210 ( .A(chng_row[10]), .ZN(n162) );
  INV_X4 U2211 ( .A(chng_row[9]), .ZN(n163) );
  INV_X4 U2212 ( .A(chng_row[8]), .ZN(n164) );
  INV_X4 U2213 ( .A(chng_row[7]), .ZN(n165) );
  INV_X4 U2214 ( .A(chng_row[6]), .ZN(n166) );
  INV_X4 U2215 ( .A(chng_row[5]), .ZN(n167) );
  INV_X4 U2216 ( .A(chng_row[4]), .ZN(n168) );
  INV_X4 U2217 ( .A(chng_row[3]), .ZN(n169) );
  INV_X4 U2218 ( .A(chng_row[2]), .ZN(n170) );
  INV_X4 U2219 ( .A(chng_row[1]), .ZN(n171) );
  INV_X4 U2220 ( .A(chng_row[0]), .ZN(n172) );
  INV_X4 U2221 ( .A(chng_col[15]), .ZN(n173) );
  INV_X4 U2222 ( .A(chng_col[14]), .ZN(n174) );
  INV_X4 U2223 ( .A(chng_col[13]), .ZN(n175) );
  INV_X4 U2224 ( .A(chng_col[12]), .ZN(n176) );
  INV_X4 U2225 ( .A(chng_col[11]), .ZN(n177) );
  INV_X4 U2226 ( .A(chng_col[10]), .ZN(n178) );
  INV_X4 U2227 ( .A(chng_col[9]), .ZN(n179) );
  INV_X4 U2228 ( .A(chng_col[8]), .ZN(n180) );
  INV_X4 U2229 ( .A(chng_col[7]), .ZN(n181) );
  INV_X4 U2230 ( .A(chng_col[6]), .ZN(n182) );
  INV_X4 U2231 ( .A(chng_col[5]), .ZN(n183) );
  INV_X4 U2232 ( .A(chng_col[4]), .ZN(n184) );
  INV_X4 U2233 ( .A(chng_col[3]), .ZN(n185) );
  INV_X4 U2234 ( .A(chng_col[2]), .ZN(n186) );
  INV_X4 U2235 ( .A(chng_col[1]), .ZN(n187) );
  INV_X4 U2236 ( .A(chng_col[0]), .ZN(n188) );
  INV_X4 U2237 ( .A(ymem_data1[255]), .ZN(n189) );
  INV_X4 U2238 ( .A(ymem_data1[254]), .ZN(n190) );
  INV_X4 U2239 ( .A(ymem_data1[253]), .ZN(n191) );
  INV_X4 U2240 ( .A(ymem_data1[251]), .ZN(n192) );
  INV_X4 U2241 ( .A(ymem_data1[250]), .ZN(n193) );
  INV_X4 U2242 ( .A(ymem_data1[249]), .ZN(n194) );
  INV_X4 U2243 ( .A(ymem_data1[239]), .ZN(n195) );
  INV_X4 U2244 ( .A(ymem_data1[238]), .ZN(n196) );
  INV_X4 U2245 ( .A(ymem_data1[237]), .ZN(n197) );
  INV_X4 U2246 ( .A(ymem_data1[236]), .ZN(n198) );
  INV_X4 U2247 ( .A(ymem_data1[235]), .ZN(n199) );
  INV_X4 U2248 ( .A(ymem_data1[234]), .ZN(n200) );
  INV_X4 U2249 ( .A(ymem_data1[233]), .ZN(n201) );
  INV_X4 U2250 ( .A(ymem_data1[232]), .ZN(n202) );
  INV_X4 U2251 ( .A(ymem_data1[231]), .ZN(n203) );
  INV_X4 U2252 ( .A(ymem_data1[230]), .ZN(n204) );
  INV_X4 U2253 ( .A(ymem_data1[229]), .ZN(n205) );
  INV_X4 U2254 ( .A(ymem_data1[228]), .ZN(n206) );
  INV_X4 U2255 ( .A(ymem_data1[227]), .ZN(n207) );
  INV_X4 U2256 ( .A(ymem_data1[226]), .ZN(n208) );
  INV_X4 U2257 ( .A(ymem_data1[225]), .ZN(n209) );
  INV_X4 U2258 ( .A(ymem_data1[224]), .ZN(n210) );
  INV_X4 U2259 ( .A(ymem_data1[223]), .ZN(n211) );
  INV_X4 U2260 ( .A(ymem_data1[222]), .ZN(n212) );
  INV_X4 U2261 ( .A(ymem_data1[221]), .ZN(n213) );
  INV_X4 U2262 ( .A(ymem_data1[220]), .ZN(n214) );
  INV_X4 U2263 ( .A(ymem_data1[219]), .ZN(n215) );
  INV_X4 U2264 ( .A(ymem_data1[218]), .ZN(n216) );
  INV_X4 U2265 ( .A(ymem_data1[217]), .ZN(n217) );
  INV_X4 U2266 ( .A(ymem_data1[216]), .ZN(n218) );
  INV_X4 U2267 ( .A(ymem_data1[215]), .ZN(n219) );
  INV_X4 U2268 ( .A(ymem_data1[214]), .ZN(n220) );
  INV_X4 U2269 ( .A(ymem_data1[213]), .ZN(n221) );
  INV_X4 U2270 ( .A(ymem_data1[212]), .ZN(n222) );
  INV_X4 U2271 ( .A(ymem_data1[211]), .ZN(n223) );
  INV_X4 U2272 ( .A(ymem_data1[210]), .ZN(n224) );
  INV_X4 U2273 ( .A(ymem_data1[209]), .ZN(n225) );
  INV_X4 U2274 ( .A(ymem_data1[208]), .ZN(n226) );
  INV_X4 U2275 ( .A(ymem_data1[207]), .ZN(n227) );
  INV_X4 U2276 ( .A(ymem_data1[206]), .ZN(n228) );
  INV_X4 U2277 ( .A(ymem_data1[205]), .ZN(n229) );
  INV_X4 U2278 ( .A(ymem_data1[204]), .ZN(n230) );
  INV_X4 U2279 ( .A(ymem_data1[203]), .ZN(n231) );
  INV_X4 U2280 ( .A(ymem_data1[202]), .ZN(n232) );
  INV_X4 U2281 ( .A(ymem_data1[201]), .ZN(n233) );
  INV_X4 U2282 ( .A(ymem_data1[200]), .ZN(n234) );
  INV_X4 U2283 ( .A(ymem_data1[199]), .ZN(n235) );
  INV_X4 U2284 ( .A(ymem_data1[198]), .ZN(n236) );
  INV_X4 U2285 ( .A(ymem_data1[197]), .ZN(n237) );
  INV_X4 U2286 ( .A(ymem_data1[196]), .ZN(n238) );
  INV_X4 U2287 ( .A(ymem_data1[195]), .ZN(n239) );
  INV_X4 U2288 ( .A(ymem_data1[194]), .ZN(n240) );
  INV_X4 U2289 ( .A(ymem_data1[193]), .ZN(n241) );
  INV_X4 U2290 ( .A(ymem_data1[192]), .ZN(n242) );
  INV_X4 U2291 ( .A(ymem_data1[191]), .ZN(n243) );
  INV_X4 U2292 ( .A(ymem_data1[190]), .ZN(n244) );
  INV_X4 U2293 ( .A(ymem_data1[189]), .ZN(n245) );
  INV_X4 U2294 ( .A(ymem_data1[188]), .ZN(n246) );
  INV_X4 U2295 ( .A(ymem_data1[187]), .ZN(n247) );
  INV_X4 U2296 ( .A(ymem_data1[186]), .ZN(n248) );
  INV_X4 U2297 ( .A(ymem_data1[185]), .ZN(n249) );
  INV_X4 U2298 ( .A(ymem_data1[184]), .ZN(n250) );
  INV_X4 U2299 ( .A(ymem_data1[183]), .ZN(n251) );
  INV_X4 U2300 ( .A(ymem_data1[182]), .ZN(n252) );
  INV_X4 U2301 ( .A(ymem_data1[181]), .ZN(n253) );
  INV_X4 U2302 ( .A(ymem_data1[180]), .ZN(n254) );
  INV_X4 U2303 ( .A(ymem_data1[179]), .ZN(n255) );
  INV_X4 U2304 ( .A(ymem_data1[178]), .ZN(n256) );
  INV_X4 U2305 ( .A(ymem_data1[177]), .ZN(n257) );
  INV_X4 U2306 ( .A(ymem_data1[176]), .ZN(n258) );
  INV_X4 U2307 ( .A(ymem_data1[175]), .ZN(n259) );
  INV_X4 U2308 ( .A(ymem_data1[174]), .ZN(n260) );
  INV_X4 U2309 ( .A(ymem_data1[173]), .ZN(n261) );
  INV_X4 U2310 ( .A(ymem_data1[172]), .ZN(n262) );
  INV_X4 U2311 ( .A(ymem_data1[171]), .ZN(n263) );
  INV_X4 U2312 ( .A(ymem_data1[170]), .ZN(n264) );
  INV_X4 U2313 ( .A(ymem_data1[169]), .ZN(n265) );
  INV_X4 U2314 ( .A(ymem_data1[168]), .ZN(n266) );
  INV_X4 U2315 ( .A(ymem_data1[167]), .ZN(n267) );
  INV_X4 U2316 ( .A(ymem_data1[166]), .ZN(n268) );
  INV_X4 U2317 ( .A(ymem_data1[165]), .ZN(n269) );
  INV_X4 U2318 ( .A(ymem_data1[164]), .ZN(n270) );
  INV_X4 U2319 ( .A(ymem_data1[163]), .ZN(n271) );
  INV_X4 U2320 ( .A(ymem_data1[162]), .ZN(n272) );
  INV_X4 U2321 ( .A(ymem_data1[161]), .ZN(n273) );
  INV_X4 U2322 ( .A(ymem_data1[160]), .ZN(n274) );
  INV_X4 U2323 ( .A(ymem_data1[159]), .ZN(n275) );
  INV_X4 U2324 ( .A(ymem_data1[158]), .ZN(n276) );
  INV_X4 U2325 ( .A(ymem_data1[157]), .ZN(n277) );
  INV_X4 U2326 ( .A(ymem_data1[156]), .ZN(n278) );
  INV_X4 U2327 ( .A(ymem_data1[155]), .ZN(n279) );
  INV_X4 U2328 ( .A(ymem_data1[154]), .ZN(n280) );
  INV_X4 U2329 ( .A(ymem_data1[153]), .ZN(n281) );
  INV_X4 U2330 ( .A(ymem_data1[152]), .ZN(n282) );
  INV_X4 U2331 ( .A(ymem_data1[151]), .ZN(n283) );
  INV_X4 U2332 ( .A(ymem_data1[150]), .ZN(n284) );
  INV_X4 U2333 ( .A(ymem_data1[149]), .ZN(n285) );
  INV_X4 U2334 ( .A(ymem_data1[148]), .ZN(n286) );
  INV_X4 U2335 ( .A(ymem_data1[147]), .ZN(n287) );
  INV_X4 U2336 ( .A(ymem_data1[146]), .ZN(n288) );
  INV_X4 U2337 ( .A(ymem_data1[145]), .ZN(n289) );
  INV_X4 U2338 ( .A(ymem_data1[144]), .ZN(n290) );
  INV_X4 U2339 ( .A(ymem_data1[143]), .ZN(n291) );
  INV_X4 U2340 ( .A(ymem_data1[142]), .ZN(n292) );
  INV_X4 U2341 ( .A(ymem_data1[141]), .ZN(n293) );
  INV_X4 U2342 ( .A(ymem_data1[140]), .ZN(n294) );
  INV_X4 U2343 ( .A(ymem_data1[139]), .ZN(n295) );
  INV_X4 U2344 ( .A(ymem_data1[138]), .ZN(n296) );
  INV_X4 U2345 ( .A(ymem_data1[137]), .ZN(n297) );
  INV_X4 U2346 ( .A(ymem_data1[136]), .ZN(n298) );
  INV_X4 U2347 ( .A(ymem_data1[135]), .ZN(n299) );
  INV_X4 U2348 ( .A(ymem_data1[134]), .ZN(n300) );
  INV_X4 U2349 ( .A(ymem_data1[133]), .ZN(n301) );
  INV_X4 U2350 ( .A(ymem_data1[132]), .ZN(n302) );
  INV_X4 U2351 ( .A(ymem_data1[131]), .ZN(n303) );
  INV_X4 U2352 ( .A(ymem_data1[130]), .ZN(n304) );
  INV_X4 U2353 ( .A(ymem_data1[129]), .ZN(n305) );
  INV_X4 U2354 ( .A(ymem_data1[128]), .ZN(n306) );
  INV_X4 U2355 ( .A(ymem_data1[127]), .ZN(n307) );
  INV_X4 U2356 ( .A(ymem_data1[126]), .ZN(n308) );
  INV_X4 U2357 ( .A(ymem_data1[125]), .ZN(n309) );
  INV_X4 U2358 ( .A(ymem_data1[124]), .ZN(n310) );
  INV_X4 U2359 ( .A(ymem_data1[123]), .ZN(n311) );
  INV_X4 U2360 ( .A(ymem_data1[122]), .ZN(n312) );
  INV_X4 U2361 ( .A(ymem_data1[121]), .ZN(n313) );
  INV_X4 U2362 ( .A(ymem_data1[120]), .ZN(n314) );
  INV_X4 U2363 ( .A(ymem_data1[119]), .ZN(n315) );
  INV_X4 U2364 ( .A(ymem_data1[118]), .ZN(n316) );
  INV_X4 U2365 ( .A(ymem_data1[117]), .ZN(n317) );
  INV_X4 U2366 ( .A(ymem_data1[116]), .ZN(n318) );
  INV_X4 U2367 ( .A(ymem_data1[115]), .ZN(n319) );
  INV_X4 U2368 ( .A(ymem_data1[114]), .ZN(n320) );
  INV_X4 U2369 ( .A(ymem_data1[113]), .ZN(n321) );
  INV_X4 U2370 ( .A(ymem_data1[112]), .ZN(n322) );
  INV_X4 U2371 ( .A(ymem_data1[111]), .ZN(n323) );
  INV_X4 U2372 ( .A(ymem_data1[110]), .ZN(n324) );
  INV_X4 U2373 ( .A(ymem_data1[109]), .ZN(n325) );
  INV_X4 U2374 ( .A(ymem_data1[108]), .ZN(n326) );
  INV_X4 U2375 ( .A(ymem_data1[107]), .ZN(n327) );
  INV_X4 U2376 ( .A(ymem_data1[106]), .ZN(n328) );
  INV_X4 U2377 ( .A(ymem_data1[105]), .ZN(n329) );
  INV_X4 U2378 ( .A(ymem_data1[104]), .ZN(n330) );
  INV_X4 U2379 ( .A(ymem_data1[103]), .ZN(n331) );
  INV_X4 U2380 ( .A(ymem_data1[102]), .ZN(n332) );
  INV_X4 U2381 ( .A(ymem_data1[101]), .ZN(n333) );
  INV_X4 U2382 ( .A(ymem_data1[100]), .ZN(n334) );
  INV_X4 U2383 ( .A(ymem_data1[99]), .ZN(n335) );
  INV_X4 U2384 ( .A(ymem_data1[98]), .ZN(n336) );
  INV_X4 U2385 ( .A(ymem_data1[97]), .ZN(n337) );
  INV_X4 U2386 ( .A(ymem_data1[96]), .ZN(n338) );
  INV_X4 U2387 ( .A(ymem_data1[95]), .ZN(n339) );
  INV_X4 U2388 ( .A(ymem_data1[94]), .ZN(n340) );
  INV_X4 U2389 ( .A(ymem_data1[93]), .ZN(n341) );
  INV_X4 U2390 ( .A(ymem_data1[92]), .ZN(n342) );
  INV_X4 U2391 ( .A(ymem_data1[91]), .ZN(n343) );
  INV_X4 U2392 ( .A(ymem_data1[90]), .ZN(n344) );
  INV_X4 U2393 ( .A(ymem_data1[89]), .ZN(n345) );
  INV_X4 U2394 ( .A(ymem_data1[88]), .ZN(n346) );
  INV_X4 U2395 ( .A(ymem_data1[87]), .ZN(n347) );
  INV_X4 U2396 ( .A(ymem_data1[86]), .ZN(n348) );
  INV_X4 U2397 ( .A(ymem_data1[85]), .ZN(n349) );
  INV_X4 U2398 ( .A(ymem_data1[84]), .ZN(n350) );
  INV_X4 U2399 ( .A(ymem_data1[83]), .ZN(n351) );
  INV_X4 U2400 ( .A(ymem_data1[82]), .ZN(n352) );
  INV_X4 U2401 ( .A(ymem_data1[81]), .ZN(n353) );
  INV_X4 U2402 ( .A(ymem_data1[80]), .ZN(n354) );
  INV_X4 U2403 ( .A(ymem_data1[79]), .ZN(n355) );
  INV_X4 U2404 ( .A(ymem_data1[78]), .ZN(n356) );
  INV_X4 U2405 ( .A(ymem_data1[77]), .ZN(n357) );
  INV_X4 U2406 ( .A(ymem_data1[76]), .ZN(n358) );
  INV_X4 U2407 ( .A(ymem_data1[75]), .ZN(n359) );
  INV_X4 U2408 ( .A(ymem_data1[74]), .ZN(n360) );
  INV_X4 U2409 ( .A(ymem_data1[73]), .ZN(n361) );
  INV_X4 U2410 ( .A(ymem_data1[72]), .ZN(n362) );
  INV_X4 U2411 ( .A(ymem_data1[71]), .ZN(n363) );
  INV_X4 U2412 ( .A(ymem_data1[70]), .ZN(n364) );
  INV_X4 U2413 ( .A(ymem_data1[69]), .ZN(n365) );
  INV_X4 U2414 ( .A(ymem_data1[68]), .ZN(n366) );
  INV_X4 U2415 ( .A(ymem_data1[67]), .ZN(n367) );
  INV_X4 U2416 ( .A(ymem_data1[66]), .ZN(n368) );
  INV_X4 U2417 ( .A(ymem_data1[65]), .ZN(n369) );
  INV_X4 U2418 ( .A(ymem_data1[64]), .ZN(n370) );
  INV_X4 U2419 ( .A(ymem_data1[63]), .ZN(n371) );
  INV_X4 U2420 ( .A(ymem_data1[62]), .ZN(n372) );
  INV_X4 U2421 ( .A(ymem_data1[61]), .ZN(n373) );
  INV_X4 U2422 ( .A(ymem_data1[60]), .ZN(n374) );
  INV_X4 U2423 ( .A(ymem_data1[59]), .ZN(n375) );
  INV_X4 U2424 ( .A(ymem_data1[58]), .ZN(n376) );
  INV_X4 U2425 ( .A(ymem_data1[57]), .ZN(n377) );
  INV_X4 U2426 ( .A(ymem_data1[56]), .ZN(n378) );
  INV_X4 U2427 ( .A(ymem_data1[55]), .ZN(n379) );
  INV_X4 U2428 ( .A(ymem_data1[54]), .ZN(n380) );
  INV_X4 U2429 ( .A(ymem_data1[53]), .ZN(n381) );
  INV_X4 U2430 ( .A(ymem_data1[52]), .ZN(n382) );
  INV_X4 U2431 ( .A(ymem_data1[51]), .ZN(n383) );
  INV_X4 U2432 ( .A(ymem_data1[50]), .ZN(n384) );
  INV_X4 U2433 ( .A(ymem_data1[49]), .ZN(n385) );
  INV_X4 U2434 ( .A(ymem_data1[48]), .ZN(n386) );
  INV_X4 U2435 ( .A(ymem_data1[47]), .ZN(n387) );
  INV_X4 U2436 ( .A(ymem_data1[46]), .ZN(n388) );
  INV_X4 U2437 ( .A(ymem_data1[45]), .ZN(n389) );
  INV_X4 U2438 ( .A(ymem_data1[44]), .ZN(n390) );
  INV_X4 U2439 ( .A(ymem_data1[43]), .ZN(n391) );
  INV_X4 U2440 ( .A(ymem_data1[42]), .ZN(n392) );
  INV_X4 U2441 ( .A(ymem_data1[41]), .ZN(n393) );
  INV_X4 U2442 ( .A(ymem_data1[40]), .ZN(n394) );
  INV_X4 U2443 ( .A(ymem_data1[39]), .ZN(n395) );
  INV_X4 U2444 ( .A(ymem_data1[38]), .ZN(n396) );
  INV_X4 U2445 ( .A(ymem_data1[37]), .ZN(n397) );
  INV_X4 U2446 ( .A(ymem_data1[36]), .ZN(n398) );
  INV_X4 U2447 ( .A(ymem_data1[35]), .ZN(n399) );
  INV_X4 U2448 ( .A(ymem_data1[34]), .ZN(n400) );
  INV_X4 U2449 ( .A(ymem_data1[33]), .ZN(n401) );
  INV_X4 U2450 ( .A(ymem_data1[32]), .ZN(n402) );
  INV_X4 U2451 ( .A(ymem_data1[31]), .ZN(n403) );
  INV_X4 U2452 ( .A(ymem_data1[30]), .ZN(n404) );
  INV_X4 U2453 ( .A(ymem_data1[29]), .ZN(n405) );
  INV_X4 U2454 ( .A(ymem_data1[28]), .ZN(n406) );
  INV_X4 U2455 ( .A(ymem_data1[27]), .ZN(n407) );
  INV_X4 U2456 ( .A(ymem_data1[26]), .ZN(n408) );
  INV_X4 U2457 ( .A(ymem_data1[25]), .ZN(n409) );
  INV_X4 U2458 ( .A(ymem_data1[24]), .ZN(n410) );
  INV_X4 U2459 ( .A(ymem_data1[23]), .ZN(n411) );
  INV_X4 U2460 ( .A(ymem_data1[22]), .ZN(n412) );
  INV_X4 U2461 ( .A(ymem_data1[21]), .ZN(n413) );
  INV_X4 U2462 ( .A(ymem_data1[20]), .ZN(n414) );
  INV_X4 U2463 ( .A(ymem_data1[19]), .ZN(n415) );
  INV_X4 U2464 ( .A(ymem_data1[18]), .ZN(n416) );
  INV_X4 U2465 ( .A(ymem_data1[17]), .ZN(n417) );
  INV_X4 U2466 ( .A(ymem_data1[16]), .ZN(n418) );
  INV_X4 U2467 ( .A(ymem_data1[15]), .ZN(n419) );
  INV_X4 U2468 ( .A(ymem_data1[14]), .ZN(n420) );
  INV_X4 U2469 ( .A(ymem_data1[13]), .ZN(n421) );
  INV_X4 U2470 ( .A(ymem_data1[12]), .ZN(n422) );
  INV_X4 U2471 ( .A(ymem_data1[11]), .ZN(n423) );
  INV_X4 U2472 ( .A(ymem_data1[10]), .ZN(n424) );
  INV_X4 U2473 ( .A(ymem_data1[9]), .ZN(n425) );
  INV_X4 U2474 ( .A(ymem_data1[8]), .ZN(n426) );
  INV_X4 U2475 ( .A(ymem_data1[7]), .ZN(n427) );
  INV_X4 U2476 ( .A(ymem_data1[6]), .ZN(n428) );
  INV_X4 U2477 ( .A(ymem_data1[5]), .ZN(n429) );
  INV_X4 U2478 ( .A(ymem_data1[4]), .ZN(n430) );
  INV_X4 U2479 ( .A(ymem_data1[3]), .ZN(n431) );
  INV_X4 U2480 ( .A(ymem_data1[2]), .ZN(n432) );
  INV_X4 U2481 ( .A(ymem_data1[1]), .ZN(n433) );
  INV_X4 U2482 ( .A(ymem_data1[0]), .ZN(n434) );
  INV_X4 U2483 ( .A(ymem_data2[255]), .ZN(n435) );
  INV_X4 U2484 ( .A(ymem_data2[254]), .ZN(n436) );
  INV_X4 U2485 ( .A(ymem_data2[253]), .ZN(n437) );
  INV_X4 U2486 ( .A(ymem_data2[252]), .ZN(n438) );
  INV_X4 U2487 ( .A(ymem_data2[251]), .ZN(n439) );
  INV_X4 U2488 ( .A(ymem_data2[250]), .ZN(n440) );
  INV_X4 U2489 ( .A(ymem_data2[249]), .ZN(n441) );
  INV_X4 U2490 ( .A(ymem_data2[248]), .ZN(n442) );
  INV_X4 U2491 ( .A(ymem_data2[247]), .ZN(n443) );
  INV_X4 U2492 ( .A(ymem_data2[246]), .ZN(n444) );
  INV_X4 U2493 ( .A(ymem_data2[245]), .ZN(n445) );
  INV_X4 U2494 ( .A(ymem_data2[244]), .ZN(n446) );
  INV_X4 U2495 ( .A(ymem_data2[243]), .ZN(n447) );
  INV_X4 U2496 ( .A(ymem_data2[242]), .ZN(n448) );
  INV_X4 U2497 ( .A(ymem_data2[241]), .ZN(n449) );
  INV_X4 U2498 ( .A(ymem_data2[240]), .ZN(n450) );
  INV_X4 U2499 ( .A(ymem_data2[175]), .ZN(n451) );
  INV_X4 U2500 ( .A(ymem_data2[174]), .ZN(n452) );
  INV_X4 U2501 ( .A(ymem_data2[173]), .ZN(n453) );
  INV_X4 U2502 ( .A(ymem_data2[172]), .ZN(n454) );
  INV_X4 U2503 ( .A(ymem_data2[171]), .ZN(n455) );
  INV_X4 U2504 ( .A(ymem_data2[170]), .ZN(n456) );
  INV_X4 U2505 ( .A(ymem_data2[169]), .ZN(n457) );
  INV_X4 U2506 ( .A(ymem_data2[168]), .ZN(n458) );
  INV_X4 U2507 ( .A(ymem_data2[167]), .ZN(n459) );
  INV_X4 U2508 ( .A(ymem_data2[166]), .ZN(n460) );
  INV_X4 U2509 ( .A(ymem_data2[165]), .ZN(n461) );
  INV_X4 U2510 ( .A(ymem_data2[164]), .ZN(n462) );
  INV_X4 U2511 ( .A(ymem_data2[163]), .ZN(n463) );
  INV_X4 U2512 ( .A(ymem_data2[162]), .ZN(n464) );
  INV_X4 U2513 ( .A(ymem_data2[161]), .ZN(n465) );
  INV_X4 U2514 ( .A(ymem_data2[160]), .ZN(n466) );
  INV_X4 U2515 ( .A(ymem_data2[159]), .ZN(n467) );
  INV_X4 U2516 ( .A(ymem_data2[158]), .ZN(n468) );
  INV_X4 U2517 ( .A(ymem_data2[157]), .ZN(n469) );
  INV_X4 U2518 ( .A(ymem_data2[156]), .ZN(n470) );
  INV_X4 U2519 ( .A(ymem_data2[155]), .ZN(n471) );
  INV_X4 U2520 ( .A(ymem_data2[154]), .ZN(n472) );
  INV_X4 U2521 ( .A(ymem_data2[153]), .ZN(n473) );
  INV_X4 U2522 ( .A(ymem_data2[152]), .ZN(n474) );
  INV_X4 U2523 ( .A(ymem_data2[151]), .ZN(n475) );
  INV_X4 U2524 ( .A(ymem_data2[150]), .ZN(n476) );
  INV_X4 U2525 ( .A(ymem_data2[149]), .ZN(n477) );
  INV_X4 U2526 ( .A(ymem_data2[148]), .ZN(n478) );
  INV_X4 U2527 ( .A(ymem_data2[147]), .ZN(n479) );
  INV_X4 U2528 ( .A(ymem_data2[146]), .ZN(n480) );
  INV_X4 U2529 ( .A(ymem_data2[145]), .ZN(n481) );
  INV_X4 U2530 ( .A(ymem_data2[144]), .ZN(n482) );
  INV_X4 U2531 ( .A(ymem_data2[143]), .ZN(n483) );
  INV_X4 U2532 ( .A(ymem_data2[142]), .ZN(n484) );
  INV_X4 U2533 ( .A(ymem_data2[141]), .ZN(n485) );
  INV_X4 U2534 ( .A(ymem_data2[140]), .ZN(n486) );
  INV_X4 U2535 ( .A(ymem_data2[139]), .ZN(n487) );
  INV_X4 U2536 ( .A(ymem_data2[138]), .ZN(n488) );
  INV_X4 U2537 ( .A(ymem_data2[137]), .ZN(n489) );
  INV_X4 U2538 ( .A(ymem_data2[136]), .ZN(n490) );
  INV_X4 U2539 ( .A(ymem_data2[135]), .ZN(n491) );
  INV_X4 U2540 ( .A(ymem_data2[134]), .ZN(n492) );
  INV_X4 U2541 ( .A(ymem_data2[133]), .ZN(n493) );
  INV_X4 U2542 ( .A(ymem_data2[132]), .ZN(n494) );
  INV_X4 U2543 ( .A(ymem_data2[131]), .ZN(n495) );
  INV_X4 U2544 ( .A(ymem_data2[130]), .ZN(n496) );
  INV_X4 U2545 ( .A(ymem_data2[129]), .ZN(n497) );
  INV_X4 U2546 ( .A(ymem_data2[128]), .ZN(n498) );
  INV_X4 U2547 ( .A(ymem_data2[127]), .ZN(n499) );
  INV_X4 U2548 ( .A(ymem_data2[126]), .ZN(n500) );
  INV_X4 U2549 ( .A(ymem_data2[125]), .ZN(n501) );
  INV_X4 U2550 ( .A(ymem_data2[124]), .ZN(n502) );
  INV_X4 U2551 ( .A(ymem_data2[123]), .ZN(n503) );
  INV_X4 U2552 ( .A(ymem_data2[122]), .ZN(n504) );
  INV_X4 U2553 ( .A(ymem_data2[121]), .ZN(n505) );
  INV_X4 U2554 ( .A(ymem_data2[120]), .ZN(n506) );
  INV_X4 U2555 ( .A(ymem_data2[119]), .ZN(n507) );
  INV_X4 U2556 ( .A(ymem_data2[118]), .ZN(n508) );
  INV_X4 U2557 ( .A(ymem_data2[117]), .ZN(n509) );
  INV_X4 U2558 ( .A(ymem_data2[116]), .ZN(n510) );
  INV_X4 U2559 ( .A(ymem_data2[115]), .ZN(n511) );
  INV_X4 U2560 ( .A(ymem_data2[114]), .ZN(n512) );
  INV_X4 U2561 ( .A(ymem_data2[113]), .ZN(n513) );
  INV_X4 U2562 ( .A(ymem_data2[112]), .ZN(n514) );
  INV_X4 U2563 ( .A(ymem_data2[111]), .ZN(n515) );
  INV_X4 U2564 ( .A(ymem_data2[110]), .ZN(n516) );
  INV_X4 U2565 ( .A(ymem_data2[109]), .ZN(n517) );
  INV_X4 U2566 ( .A(ymem_data2[108]), .ZN(n518) );
  INV_X4 U2567 ( .A(ymem_data2[107]), .ZN(n519) );
  INV_X4 U2568 ( .A(ymem_data2[106]), .ZN(n520) );
  INV_X4 U2569 ( .A(ymem_data2[105]), .ZN(n521) );
  INV_X4 U2570 ( .A(ymem_data2[104]), .ZN(n522) );
  INV_X4 U2571 ( .A(ymem_data2[103]), .ZN(n523) );
  INV_X4 U2572 ( .A(ymem_data2[102]), .ZN(n524) );
  INV_X4 U2573 ( .A(ymem_data2[101]), .ZN(n525) );
  INV_X4 U2574 ( .A(ymem_data2[100]), .ZN(n526) );
  INV_X4 U2575 ( .A(ymem_data2[99]), .ZN(n527) );
  INV_X4 U2576 ( .A(ymem_data2[98]), .ZN(n528) );
  INV_X4 U2577 ( .A(ymem_data2[97]), .ZN(n529) );
  INV_X4 U2578 ( .A(ymem_data2[96]), .ZN(n530) );
  INV_X4 U2579 ( .A(ymem_data2[95]), .ZN(n531) );
  INV_X4 U2580 ( .A(ymem_data2[94]), .ZN(n532) );
  INV_X4 U2581 ( .A(ymem_data2[93]), .ZN(n533) );
  INV_X4 U2582 ( .A(ymem_data2[92]), .ZN(n534) );
  INV_X4 U2583 ( .A(ymem_data2[91]), .ZN(n535) );
  INV_X4 U2584 ( .A(ymem_data2[90]), .ZN(n536) );
  INV_X4 U2585 ( .A(ymem_data2[89]), .ZN(n537) );
  INV_X4 U2586 ( .A(ymem_data2[88]), .ZN(n538) );
  INV_X4 U2587 ( .A(ymem_data2[87]), .ZN(n539) );
  INV_X4 U2588 ( .A(ymem_data2[86]), .ZN(n540) );
  INV_X4 U2589 ( .A(ymem_data2[85]), .ZN(n541) );
  INV_X4 U2590 ( .A(ymem_data2[84]), .ZN(n542) );
  INV_X4 U2591 ( .A(ymem_data2[83]), .ZN(n543) );
  INV_X4 U2592 ( .A(ymem_data2[82]), .ZN(n544) );
  INV_X4 U2593 ( .A(ymem_data2[81]), .ZN(n545) );
  INV_X4 U2594 ( .A(ymem_data2[80]), .ZN(n546) );
  INV_X4 U2595 ( .A(ymem_data2[79]), .ZN(n547) );
  INV_X4 U2596 ( .A(ymem_data2[78]), .ZN(n548) );
  INV_X4 U2597 ( .A(ymem_data2[77]), .ZN(n549) );
  INV_X4 U2598 ( .A(ymem_data2[76]), .ZN(n550) );
  INV_X4 U2599 ( .A(ymem_data2[75]), .ZN(n551) );
  INV_X4 U2600 ( .A(ymem_data2[74]), .ZN(n552) );
  INV_X4 U2601 ( .A(ymem_data2[73]), .ZN(n553) );
  INV_X4 U2602 ( .A(ymem_data2[72]), .ZN(n554) );
  INV_X4 U2603 ( .A(ymem_data2[71]), .ZN(n555) );
  INV_X4 U2604 ( .A(ymem_data2[70]), .ZN(n556) );
  INV_X4 U2605 ( .A(ymem_data2[69]), .ZN(n557) );
  INV_X4 U2606 ( .A(ymem_data2[68]), .ZN(n558) );
  INV_X4 U2607 ( .A(ymem_data2[67]), .ZN(n559) );
  INV_X4 U2608 ( .A(ymem_data2[66]), .ZN(n560) );
  INV_X4 U2609 ( .A(ymem_data2[65]), .ZN(n561) );
  INV_X4 U2610 ( .A(ymem_data2[64]), .ZN(n562) );
  INV_X4 U2611 ( .A(ymem_data2[63]), .ZN(n563) );
  INV_X4 U2612 ( .A(ymem_data2[62]), .ZN(n564) );
  INV_X4 U2613 ( .A(ymem_data2[61]), .ZN(n565) );
  INV_X4 U2614 ( .A(ymem_data2[60]), .ZN(n566) );
  INV_X4 U2615 ( .A(ymem_data2[59]), .ZN(n567) );
  INV_X4 U2616 ( .A(ymem_data2[58]), .ZN(n568) );
  INV_X4 U2617 ( .A(ymem_data2[57]), .ZN(n569) );
  INV_X4 U2618 ( .A(ymem_data2[56]), .ZN(n570) );
  INV_X4 U2619 ( .A(ymem_data2[55]), .ZN(n571) );
  INV_X4 U2620 ( .A(ymem_data2[54]), .ZN(n572) );
  INV_X4 U2621 ( .A(ymem_data2[53]), .ZN(n573) );
  INV_X4 U2622 ( .A(ymem_data2[52]), .ZN(n574) );
  INV_X4 U2623 ( .A(ymem_data2[51]), .ZN(n575) );
  INV_X4 U2624 ( .A(ymem_data2[50]), .ZN(n576) );
  INV_X4 U2625 ( .A(ymem_data2[49]), .ZN(n577) );
  INV_X4 U2626 ( .A(ymem_data2[48]), .ZN(n578) );
  INV_X4 U2627 ( .A(ymem_data2[47]), .ZN(n579) );
  INV_X4 U2628 ( .A(ymem_data2[46]), .ZN(n580) );
  INV_X4 U2629 ( .A(ymem_data2[45]), .ZN(n581) );
  INV_X4 U2630 ( .A(ymem_data2[44]), .ZN(n582) );
  INV_X4 U2631 ( .A(ymem_data2[43]), .ZN(n583) );
  INV_X4 U2632 ( .A(ymem_data2[42]), .ZN(n584) );
  INV_X4 U2633 ( .A(ymem_data2[41]), .ZN(n585) );
  INV_X4 U2634 ( .A(ymem_data2[40]), .ZN(n586) );
  INV_X4 U2635 ( .A(ymem_data2[39]), .ZN(n587) );
  INV_X4 U2636 ( .A(ymem_data2[38]), .ZN(n588) );
  INV_X4 U2637 ( .A(ymem_data2[37]), .ZN(n589) );
  INV_X4 U2638 ( .A(ymem_data2[36]), .ZN(n590) );
  INV_X4 U2639 ( .A(ymem_data2[35]), .ZN(n591) );
  INV_X4 U2640 ( .A(ymem_data2[34]), .ZN(n592) );
  INV_X4 U2641 ( .A(ymem_data2[33]), .ZN(n593) );
  INV_X4 U2642 ( .A(ymem_data2[32]), .ZN(n594) );
  INV_X4 U2643 ( .A(ymem_data2[31]), .ZN(n595) );
  INV_X4 U2644 ( .A(ymem_data2[30]), .ZN(n596) );
  INV_X4 U2645 ( .A(ymem_data2[29]), .ZN(n597) );
  INV_X4 U2646 ( .A(ymem_data2[28]), .ZN(n598) );
  INV_X4 U2647 ( .A(ymem_data2[27]), .ZN(n599) );
  INV_X4 U2648 ( .A(ymem_data2[26]), .ZN(n600) );
  INV_X4 U2649 ( .A(ymem_data2[25]), .ZN(n601) );
  INV_X4 U2650 ( .A(ymem_data2[24]), .ZN(n602) );
  INV_X4 U2651 ( .A(ymem_data2[23]), .ZN(n603) );
  INV_X4 U2652 ( .A(ymem_data2[22]), .ZN(n604) );
  INV_X4 U2653 ( .A(ymem_data2[21]), .ZN(n605) );
  INV_X4 U2654 ( .A(ymem_data2[20]), .ZN(n606) );
  INV_X4 U2655 ( .A(ymem_data2[19]), .ZN(n607) );
  INV_X4 U2656 ( .A(ymem_data2[18]), .ZN(n608) );
  INV_X4 U2657 ( .A(ymem_data2[17]), .ZN(n609) );
  INV_X4 U2658 ( .A(ymem_data2[16]), .ZN(n610) );
  INV_X4 U2659 ( .A(ymem_data2[15]), .ZN(n611) );
  INV_X4 U2660 ( .A(ymem_data2[14]), .ZN(n612) );
  INV_X4 U2661 ( .A(ymem_data2[13]), .ZN(n613) );
  INV_X4 U2662 ( .A(ymem_data2[12]), .ZN(n614) );
  INV_X4 U2663 ( .A(ymem_data2[11]), .ZN(n615) );
  INV_X4 U2664 ( .A(ymem_data2[10]), .ZN(n616) );
  INV_X4 U2665 ( .A(ymem_data2[9]), .ZN(n617) );
  INV_X4 U2666 ( .A(ymem_data2[8]), .ZN(n618) );
  INV_X4 U2667 ( .A(ymem_data2[7]), .ZN(n619) );
  INV_X4 U2668 ( .A(ymem_data2[6]), .ZN(n620) );
  INV_X4 U2669 ( .A(ymem_data2[5]), .ZN(n621) );
  INV_X4 U2670 ( .A(ymem_data2[4]), .ZN(n622) );
  INV_X4 U2671 ( .A(ymem_data2[3]), .ZN(n623) );
  INV_X4 U2672 ( .A(ymem_data2[2]), .ZN(n624) );
  INV_X4 U2673 ( .A(ymem_data2[1]), .ZN(n625) );
  INV_X4 U2674 ( .A(ymem_data2[0]), .ZN(n626) );
  OR3_X1 U2675 ( .A1(n751), .A2(n100), .A3(n752), .ZN(n713) );
  AND2_X1 U2676 ( .A1(n3277), .A2(n9), .ZN(n718) );
  AND2_X1 U2677 ( .A1(n109), .A2(n728), .ZN(n699) );
  AND2_X1 U2679 ( .A1(n3309), .A2(reset), .ZN(n1753) );
  AND2_X1 U2681 ( .A1(n118), .A2(n1778), .ZN(n799) );
  AND2_X1 U2682 ( .A1(n3271), .A2(n9), .ZN(n813) );
  AND2_X1 U2683 ( .A1(n3261), .A2(n9), .ZN(n805) );
  AND2_X1 U2685 ( .A1(chng_img[9]), .A2(n3204), .ZN(U93_Z_9) );
  AND2_X1 U2686 ( .A1(chng_img[8]), .A2(n3204), .ZN(U93_Z_8) );
  AND2_X1 U2687 ( .A1(chng_img[7]), .A2(n3204), .ZN(U93_Z_7) );
  AND2_X1 U2688 ( .A1(chng_img[6]), .A2(n3204), .ZN(U93_Z_6) );
  AND2_X1 U2689 ( .A1(chng_img[5]), .A2(n3204), .ZN(U93_Z_5) );
  AND2_X1 U2690 ( .A1(chng_real[23]), .A2(n3204), .ZN(U93_Z_47) );
  AND2_X1 U2691 ( .A1(chng_real[22]), .A2(n3204), .ZN(U93_Z_46) );
  AND2_X1 U2692 ( .A1(chng_real[21]), .A2(n3204), .ZN(U93_Z_45) );
  AND2_X1 U2693 ( .A1(chng_real[20]), .A2(n3204), .ZN(U93_Z_44) );
  AND2_X1 U2694 ( .A1(chng_real[19]), .A2(n3204), .ZN(U93_Z_43) );
  AND2_X1 U2695 ( .A1(chng_real[18]), .A2(n3204), .ZN(U93_Z_42) );
  AND2_X1 U2696 ( .A1(chng_real[17]), .A2(n3204), .ZN(U93_Z_41) );
  AND2_X1 U2697 ( .A1(chng_real[16]), .A2(n3204), .ZN(U93_Z_40) );
  AND2_X1 U2698 ( .A1(chng_img[4]), .A2(n3204), .ZN(U93_Z_4) );
  AND2_X1 U2699 ( .A1(chng_real[15]), .A2(n3204), .ZN(U93_Z_39) );
  AND2_X1 U2700 ( .A1(chng_real[14]), .A2(n3204), .ZN(U93_Z_38) );
  AND2_X1 U2701 ( .A1(chng_real[13]), .A2(n3204), .ZN(U93_Z_37) );
  AND2_X1 U2702 ( .A1(chng_real[12]), .A2(n3204), .ZN(U93_Z_36) );
  AND2_X1 U2703 ( .A1(chng_real[11]), .A2(n3204), .ZN(U93_Z_35) );
  AND2_X1 U2704 ( .A1(chng_real[10]), .A2(n3204), .ZN(U93_Z_34) );
  AND2_X1 U2705 ( .A1(chng_real[9]), .A2(n3204), .ZN(U93_Z_33) );
  AND2_X1 U2706 ( .A1(chng_real[8]), .A2(n3204), .ZN(U93_Z_32) );
  AND2_X1 U2707 ( .A1(chng_real[7]), .A2(n3204), .ZN(U93_Z_31) );
  AND2_X1 U2708 ( .A1(chng_real[6]), .A2(n3204), .ZN(U93_Z_30) );
  AND2_X1 U2709 ( .A1(chng_img[3]), .A2(n3204), .ZN(U93_Z_3) );
  AND2_X1 U2710 ( .A1(chng_real[5]), .A2(n3204), .ZN(U93_Z_29) );
  AND2_X1 U2711 ( .A1(chng_real[4]), .A2(n3204), .ZN(U93_Z_28) );
  AND2_X1 U2712 ( .A1(chng_real[3]), .A2(n3204), .ZN(U93_Z_27) );
  AND2_X1 U2713 ( .A1(chng_real[2]), .A2(n3204), .ZN(U93_Z_26) );
  AND2_X1 U2714 ( .A1(chng_real[1]), .A2(n3204), .ZN(U93_Z_25) );
  AND2_X1 U2715 ( .A1(chng_real[0]), .A2(n3204), .ZN(U93_Z_24) );
  AND2_X1 U2716 ( .A1(chng_img[23]), .A2(n3204), .ZN(U93_Z_23) );
  AND2_X1 U2717 ( .A1(chng_img[22]), .A2(n3204), .ZN(U93_Z_22) );
  AND2_X1 U2718 ( .A1(chng_img[21]), .A2(n3204), .ZN(U93_Z_21) );
  AND2_X1 U2719 ( .A1(chng_img[20]), .A2(n3204), .ZN(U93_Z_20) );
  AND2_X1 U2720 ( .A1(chng_img[2]), .A2(n3204), .ZN(U93_Z_2) );
  AND2_X1 U2721 ( .A1(chng_img[19]), .A2(n3204), .ZN(U93_Z_19) );
  AND2_X1 U2722 ( .A1(chng_img[18]), .A2(n3204), .ZN(U93_Z_18) );
  AND2_X1 U2723 ( .A1(chng_img[17]), .A2(n3204), .ZN(U93_Z_17) );
  AND2_X1 U2724 ( .A1(chng_img[16]), .A2(n3204), .ZN(U93_Z_16) );
  AND2_X1 U2725 ( .A1(chng_img[15]), .A2(n3204), .ZN(U93_Z_15) );
  AND2_X1 U2726 ( .A1(chng_img[14]), .A2(n3204), .ZN(U93_Z_14) );
  AND2_X1 U2727 ( .A1(chng_img[13]), .A2(n3204), .ZN(U93_Z_13) );
  AND2_X1 U2728 ( .A1(chng_img[12]), .A2(n3204), .ZN(U93_Z_12) );
  AND2_X1 U2729 ( .A1(chng_img[11]), .A2(n3204), .ZN(U93_Z_11) );
  AND2_X1 U2730 ( .A1(chng_img[10]), .A2(n3204), .ZN(U93_Z_10) );
  AND2_X1 U2731 ( .A1(chng_img[1]), .A2(n3204), .ZN(U93_Z_1) );
  AND2_X1 U2732 ( .A1(chng_img[0]), .A2(n3204), .ZN(U93_Z_0) );
  AND2_X1 U2734 ( .A1(n2146), .A2(n825), .ZN(n1778) );
  AND2_X1 U2737 ( .A1(n2503), .A2(n3257), .ZN(n693) );
  AND2_X1 U2739 ( .A1(n2506), .A2(n2503), .ZN(n732) );
  OR4_X1 U2740 ( .A1(n2529), .A2(n2553), .A3(n2554), .A4(n2555), .ZN(n2552) );
  OR4_X1 U2741 ( .A1(n2556), .A2(n2547), .A3(n2546), .A4(n2557), .ZN(n2551) );
  DFF_X2 current_state_reg_1_ ( .D(U95_Z_1), .CK(clock), .Q(n[2371]), .QN(n151) );
  DFF_X2 current_state_reg_0_ ( .D(U95_Z_0), .CK(clock), .Q(n[2370]), .QN(n152) );
  DFF_X2 current_state_reg_2_ ( .D(U95_Z_2), .CK(clock), .Q(n[2372]), .QN(n149) );
  DFF_X2 temp_yVal_reg_47_ ( .D(n2678), .CK(clock), .Q(U72_DATA1_47), .QN(n11)
         );
  DFF_X2 temp_yVal_reg_46_ ( .D(n2677), .CK(clock), .Q(U72_DATA1_46), .QN(n12)
         );
  DFF_X2 temp_yVal_reg_45_ ( .D(n2676), .CK(clock), .Q(U72_DATA1_45), .QN(n13)
         );
  DFF_X2 temp_yVal_reg_44_ ( .D(n2675), .CK(clock), .Q(U72_DATA1_44), .QN(n14)
         );
  DFF_X2 temp_yVal_reg_43_ ( .D(n2674), .CK(clock), .Q(U72_DATA1_43), .QN(n15)
         );
  DFF_X2 temp_yVal_reg_42_ ( .D(n2673), .CK(clock), .Q(U72_DATA1_42), .QN(n16)
         );
  DFF_X2 temp_yVal_reg_41_ ( .D(n2672), .CK(clock), .Q(U72_DATA1_41), .QN(n17)
         );
  DFF_X2 temp_yVal_reg_40_ ( .D(n2671), .CK(clock), .Q(U72_DATA1_40), .QN(n18)
         );
  DFF_X2 temp_yVal_reg_39_ ( .D(n2670), .CK(clock), .Q(U72_DATA1_39), .QN(n19)
         );
  DFF_X2 temp_yVal_reg_38_ ( .D(n2669), .CK(clock), .Q(U72_DATA1_38), .QN(n20)
         );
  DFF_X2 temp_yVal_reg_37_ ( .D(n2668), .CK(clock), .Q(U72_DATA1_37), .QN(n21)
         );
  DFF_X2 temp_yVal_reg_36_ ( .D(n2667), .CK(clock), .Q(U72_DATA1_36), .QN(n22)
         );
  DFF_X2 temp_yVal_reg_35_ ( .D(n2666), .CK(clock), .Q(U72_DATA1_35), .QN(n23)
         );
  DFF_X2 temp_yVal_reg_34_ ( .D(n2665), .CK(clock), .Q(U72_DATA1_34), .QN(n24)
         );
  DFF_X2 temp_yVal_reg_33_ ( .D(n2664), .CK(clock), .Q(U72_DATA1_33), .QN(n25)
         );
  DFF_X2 temp_yVal_reg_32_ ( .D(n2663), .CK(clock), .Q(U72_DATA1_32), .QN(n26)
         );
  DFF_X2 temp_yVal_reg_31_ ( .D(n2662), .CK(clock), .Q(U72_DATA1_31), .QN(n27)
         );
  DFF_X2 temp_yVal_reg_30_ ( .D(n2661), .CK(clock), .Q(U72_DATA1_30), .QN(n28)
         );
  DFF_X2 temp_yVal_reg_29_ ( .D(n2660), .CK(clock), .Q(U72_DATA1_29), .QN(n29)
         );
  NAND3_X2 U4 ( .A1(n152), .A2(n151), .A3(n[2372]), .ZN(n829) );
  NAND2_X4 U12 ( .A1(n812), .A2(exModDone), .ZN(n3198) );
  NAND2_X4 U17 ( .A1(n1753), .A2(n130), .ZN(n3200) );
  NAND2_X4 U19 ( .A1(n1753), .A2(n3287), .ZN(n3201) );
  INV_X2 U22 ( .A(n865), .ZN(n3245) );
  OR2_X4 U24 ( .A1(n1772), .A2(n3301), .ZN(n834) );
  NOR2_X4 U27 ( .A1(n717), .A2(n156), .ZN(n3202) );
  INV_X2 U29 ( .A(n864), .ZN(n3247) );
  OR2_X4 U32 ( .A1(n2504), .A2(n146), .ZN(n3203) );
  AND2_X4 U34 ( .A1(n2153), .A2(reset), .ZN(n3204) );
  AND2_X4 U37 ( .A1(n2235), .A2(n2501), .ZN(n3205) );
  INV_X2 U39 ( .A(n866), .ZN(n3243) );
  AND2_X4 U42 ( .A1(n804), .A2(exModDone), .ZN(n3206) );
  OR2_X4 U44 ( .A1(n823), .A2(n156), .ZN(n3207) );
  OR2_X4 U47 ( .A1(n2145), .A2(n698), .ZN(n3208) );
  OR2_X4 U49 ( .A1(n814), .A2(n3258), .ZN(n3209) );
  OR2_X4 U52 ( .A1(n710), .A2(n2145), .ZN(n3210) );
  NAND2_X2 U54 ( .A1(n727), .A2(exModDone), .ZN(n3211) );
  AND2_X4 U57 ( .A1(n1753), .A2(n150), .ZN(n3212) );
  NAND2_X2 U59 ( .A1(n1753), .A2(n3291), .ZN(n3213) );
  AND2_X4 U61 ( .A1(n775), .A2(n776), .ZN(n3214) );
  AND2_X4 U63 ( .A1(n[2370]), .A2(n1798), .ZN(n3215) );
  AND2_X4 U66 ( .A1(n3278), .A2(n793), .ZN(n3216) );
  OR2_X4 U69 ( .A1(n156), .A2(n9), .ZN(n3217) );
  INV_X4 U72 ( .A(n723), .ZN(n3296) );
  INV_X4 U73 ( .A(n723), .ZN(n3297) );
  INV_X4 U74 ( .A(n3209), .ZN(n3276) );
  INV_X4 U77 ( .A(n3209), .ZN(n3277) );
  INV_X4 U78 ( .A(n3285), .ZN(n3284) );
  INV_X4 U79 ( .A(n815), .ZN(n3292) );
  INV_X4 U81 ( .A(n3245), .ZN(n3244) );
  INV_X4 U88 ( .A(n3265), .ZN(n3264) );
  INV_X4 U91 ( .A(n3243), .ZN(n3242) );
  INV_X4 U104 ( .A(n1782), .ZN(n3295) );
  INV_X4 U107 ( .A(n3247), .ZN(n3246) );
  INV_X4 U108 ( .A(n3208), .ZN(n3263) );
  INV_X4 U111 ( .A(n3210), .ZN(n3270) );
  INV_X4 U113 ( .A(n3208), .ZN(n3262) );
  INV_X4 U114 ( .A(n3210), .ZN(n3271) );
  INV_X4 U115 ( .A(n1764), .ZN(n3294) );
  INV_X4 U118 ( .A(n3239), .ZN(n3238) );
  INV_X4 U119 ( .A(n778), .ZN(n3285) );
  INV_X4 U120 ( .A(n3256), .ZN(n3255) );
  INV_X4 U123 ( .A(n3260), .ZN(n3261) );
  INV_X4 U125 ( .A(n3250), .ZN(n3248) );
  INV_X4 U128 ( .A(n3250), .ZN(n3249) );
  INV_X4 U129 ( .A(n3252), .ZN(n3251) );
  INV_X4 U132 ( .A(n3216), .ZN(n3283) );
  INV_X4 U134 ( .A(n3216), .ZN(n3282) );
  INV_X4 U137 ( .A(n3213), .ZN(n3273) );
  NOR3_X2 U139 ( .A1(n141), .A2(n121), .A3(n113), .ZN(n2418) );
  INV_X4 U143 ( .A(n851), .ZN(n3267) );
  INV_X4 U146 ( .A(n852), .ZN(n3265) );
  NAND4_X2 U147 ( .A1(n2473), .A2(n2501), .A3(n793), .A4(n791), .ZN(n2472) );
  AOI222_X1 U152 ( .A1(n145), .A2(n699), .B1(n121), .B2(n94), .C1(n141), .C2(
        n784), .ZN(n768) );
  NOR2_X2 U157 ( .A1(n3280), .A2(n113), .ZN(n2246) );
  INV_X4 U160 ( .A(n857), .ZN(n3256) );
  INV_X4 U161 ( .A(n1764), .ZN(n3293) );
  INV_X4 U164 ( .A(n3254), .ZN(n3253) );
  INV_X4 U166 ( .A(n860), .ZN(n3254) );
  INV_X4 U167 ( .A(n870), .ZN(n3239) );
  INV_X4 U177 ( .A(n862), .ZN(n3252) );
  INV_X4 U180 ( .A(n863), .ZN(n3250) );
  INV_X4 U181 ( .A(n3290), .ZN(n3289) );
  INV_X4 U184 ( .A(n628), .ZN(n3290) );
  INV_X4 U186 ( .A(n3213), .ZN(n3272) );
  INV_X4 U187 ( .A(n3212), .ZN(n3275) );
  AOI22_X2 U192 ( .A1(n115), .A2(n741), .B1(n3220), .B2(n742), .ZN(n740) );
  OAI21_X2 U197 ( .B1(n750), .B2(n713), .A(n146), .ZN(n738) );
  AOI22_X2 U200 ( .A1(n136), .A2(n703), .B1(n3220), .B2(n705), .ZN(n702) );
  OAI21_X2 U201 ( .B1(n712), .B2(n713), .A(n146), .ZN(n700) );
  OAI211_X2 U204 ( .C1(n3203), .C2(n687), .A(n688), .B(n689), .ZN(n641) );
  INV_X4 U206 ( .A(n775), .ZN(n113) );
  AOI22_X2 U207 ( .A1(n97), .A2(n3220), .B1(n751), .B2(n146), .ZN(n1765) );
  INV_X4 U212 ( .A(n3259), .ZN(n3258) );
  INV_X4 U217 ( .A(n3241), .ZN(n3240) );
  INV_X4 U220 ( .A(n869), .ZN(n3241) );
  OAI222_X2 U221 ( .A1(n791), .A2(n706), .B1(n776), .B2(n709), .C1(n792), .C2(
        n793), .ZN(n790) );
  AOI21_X2 U224 ( .B1(n745), .B2(n3280), .A(n718), .ZN(n816) );
  OAI211_X2 U226 ( .C1(n3203), .C2(n729), .A(n688), .B(n730), .ZN(n646) );
  OAI21_X2 U227 ( .B1(n131), .B2(n3), .A(reset), .ZN(n637) );
  AOI22_X2 U232 ( .A1(n146), .A2(n100), .B1(n3220), .B2(n745), .ZN(n1767) );
  AOI22_X2 U237 ( .A1(n784), .A2(n3220), .B1(n752), .B2(n146), .ZN(n1770) );
  NAND2_X2 U240 ( .A1(n2248), .A2(n2140), .ZN(n2301) );
  AOI22_X2 U241 ( .A1(n712), .A2(n146), .B1(n107), .B2(n122), .ZN(n1763) );
  AOI22_X2 U244 ( .A1(n90), .A2(n3220), .B1(n752), .B2(n146), .ZN(n1784) );
  INV_X4 U247 ( .A(n3269), .ZN(n3268) );
  INV_X4 U252 ( .A(n849), .ZN(n3269) );
  AOI22_X2 U257 ( .A1(n3220), .A2(n132), .B1(n146), .B2(n105), .ZN(n870) );
  AOI222_X1 U260 ( .A1(n146), .A2(n699), .B1(n3220), .B2(n737), .C1(n136), 
        .C2(n109), .ZN(n1764) );
  AOI222_X1 U261 ( .A1(n3220), .A2(n737), .B1(n146), .B2(n736), .C1(n115), 
        .C2(n111), .ZN(n1782) );
  INV_X4 U264 ( .A(n3233), .ZN(n3232) );
  INV_X4 U266 ( .A(n3207), .ZN(n3234) );
  INV_X4 U267 ( .A(n3207), .ZN(n3235) );
  AOI22_X2 U272 ( .A1(n750), .A2(n3279), .B1(n105), .B2(n113), .ZN(n824) );
  INV_X4 U277 ( .A(n1766), .ZN(n132) );
  AOI22_X2 U280 ( .A1(n3220), .A2(n132), .B1(n146), .B2(n112), .ZN(n862) );
  INV_X4 U281 ( .A(n3281), .ZN(n3280) );
  INV_X4 U284 ( .A(n782), .ZN(n3281) );
  INV_X4 U286 ( .A(n3279), .ZN(n3278) );
  INV_X4 U287 ( .A(n3214), .ZN(n3288) );
  INV_X4 U292 ( .A(n3212), .ZN(n3274) );
  INV_X4 U297 ( .A(n822), .ZN(n7) );
  INV_X4 U300 ( .A(n632), .ZN(n72) );
  INV_X4 U301 ( .A(reset), .ZN(n3300) );
  AOI222_X1 U304 ( .A1(n799), .A2(n117), .B1(n130), .B2(n719), .C1(n113), .C2(
        n749), .ZN(n798) );
  INV_X4 U306 ( .A(n3226), .ZN(n3227) );
  INV_X4 U307 ( .A(n3229), .ZN(n3228) );
  INV_X4 U312 ( .A(n3206), .ZN(n3231) );
  INV_X4 U317 ( .A(n2156), .ZN(n3291) );
  INV_X4 U320 ( .A(n3257), .ZN(n3259) );
  OAI222_X2 U321 ( .A1(n694), .A2(n695), .B1(n696), .B2(n3203), .C1(n697), 
        .C2(n698), .ZN(n640) );
  NOR3_X2 U324 ( .A1(n145), .A2(n141), .A3(n3287), .ZN(n2235) );
  AOI22_X2 U326 ( .A1(n751), .A2(n3282), .B1(n132), .B2(n3280), .ZN(n803) );
  AOI222_X1 U327 ( .A1(n720), .A2(n130), .B1(n752), .B2(n3282), .C1(n737), 
        .C2(n3280), .ZN(n770) );
  NOR2_X2 U332 ( .A1(n2291), .A2(n113), .ZN(n2420) );
  INV_X4 U337 ( .A(n695), .ZN(n146) );
  AOI21_X2 U340 ( .B1(n2157), .B2(n2158), .A(n3301), .ZN(U90_Z_0) );
  OAI222_X2 U341 ( .A1(n729), .A2(n795), .B1(n775), .B2(n2180), .C1(n2181), 
        .C2(n797), .ZN(n2179) );
  AOI21_X2 U344 ( .B1(n698), .B2(n708), .A(n776), .ZN(n773) );
  AOI21_X2 U346 ( .B1(n735), .B2(n746), .A(n775), .ZN(n774) );
  OAI21_X2 U347 ( .B1(n812), .B2(n813), .A(n3287), .ZN(n811) );
  INV_X4 U352 ( .A(n1807), .ZN(n3233) );
  INV_X4 U357 ( .A(n3203), .ZN(n3220) );
  INV_X4 U360 ( .A(n3222), .ZN(n3223) );
  OAI222_X2 U361 ( .A1(n696), .A2(n3203), .B1(n733), .B2(n695), .C1(n734), 
        .C2(n735), .ZN(n645) );
  NOR2_X2 U364 ( .A1(n2291), .A2(n139), .ZN(n2248) );
  NOR2_X2 U366 ( .A1(n2302), .A2(n2291), .ZN(n2419) );
  AOI22_X2 U367 ( .A1(n712), .A2(n827), .B1(n727), .B2(n765), .ZN(n826) );
  AOI21_X2 U372 ( .B1(n735), .B2(n814), .A(n3216), .ZN(n810) );
  INV_X4 U377 ( .A(n794), .ZN(n3279) );
  NOR2_X2 U380 ( .A1(n2291), .A2(n145), .ZN(n2247) );
  INV_X4 U381 ( .A(n3211), .ZN(n3225) );
  OAI21_X2 U384 ( .B1(n764), .B2(n765), .A(reset), .ZN(n632) );
  OAI21_X2 U386 ( .B1(n764), .B2(n828), .A(reset), .ZN(n822) );
  INV_X4 U387 ( .A(n3217), .ZN(n3237) );
  INV_X4 U392 ( .A(n3217), .ZN(n3236) );
  OAI22_X2 U397 ( .A1(n714), .A2(n3286), .B1(n716), .B2(n717), .ZN(n643) );
  NAND2_X2 U400 ( .A1(n717), .A2(n3286), .ZN(n765) );
  INV_X4 U401 ( .A(n634), .ZN(n150) );
  INV_X4 U404 ( .A(n717), .ZN(n130) );
  INV_X4 U406 ( .A(n1810), .ZN(n3229) );
  INV_X4 U407 ( .A(n3206), .ZN(n3230) );
  INV_X4 U412 ( .A(n856), .ZN(n3257) );
  OAI21_X2 U417 ( .B1(n724), .B2(n715), .A(n725), .ZN(n642) );
  OAI21_X2 U420 ( .B1(n726), .B2(n727), .A(n130), .ZN(n725) );
  AOI21_X2 U421 ( .B1(n728), .B2(n698), .A(n722), .ZN(n726) );
  OAI21_X2 U424 ( .B1(n3301), .B2(n1785), .A(n134), .ZN(U95_Z_2) );
  OAI21_X2 U426 ( .B1(n3236), .B2(n1788), .A(n3287), .ZN(n1786) );
  AOI21_X2 U427 ( .B1(n724), .B2(n714), .A(n156), .ZN(n1788) );
  INV_X4 U432 ( .A(n3211), .ZN(n3224) );
  INV_X4 U437 ( .A(reset), .ZN(n3301) );
  NOR3_X2 U440 ( .A1(n2153), .A2(n765), .A3(n2155), .ZN(n2154) );
  OAI211_X2 U441 ( .C1(n1799), .C2(n829), .A(reset), .B(n831), .ZN(n2155) );
  AOI222_X1 U444 ( .A1(ymem_data1[114]), .A2(n150), .B1(ymem_data1[242]), .B2(
        n765), .C1(ymem_data1[50]), .C2(n3291), .ZN(n2519) );
  AOI222_X1 U446 ( .A1(ymem_data1[113]), .A2(n150), .B1(ymem_data1[241]), .B2(
        n765), .C1(ymem_data1[49]), .C2(n3291), .ZN(n2527) );
  AOI222_X1 U447 ( .A1(ymem_data1[117]), .A2(n150), .B1(ymem_data1[245]), .B2(
        n765), .C1(ymem_data1[53]), .C2(n3291), .ZN(n2538) );
  AOI222_X1 U452 ( .A1(ymem_data1[118]), .A2(n150), .B1(ymem_data1[246]), .B2(
        n765), .C1(ymem_data1[54]), .C2(n3291), .ZN(n2541) );
  AOI211_X2 U457 ( .C1(ymem_data2[46]), .C2(n3242), .A(n1743), .B(n1744), .ZN(
        n1727) );
  AOI211_X2 U460 ( .C1(n3272), .C2(n1729), .A(n1730), .B(n1731), .ZN(n1728) );
  AOI211_X2 U461 ( .C1(ymem_data2[45]), .C2(n3242), .A(n1724), .B(n1725), .ZN(
        n1708) );
  AOI211_X2 U464 ( .C1(n3272), .C2(n1710), .A(n1711), .B(n1712), .ZN(n1709) );
  AOI211_X2 U466 ( .C1(ymem_data2[44]), .C2(n866), .A(n1705), .B(n1706), .ZN(
        n1689) );
  AOI211_X2 U467 ( .C1(n3272), .C2(n1691), .A(n1692), .B(n1693), .ZN(n1690) );
  AOI211_X2 U472 ( .C1(ymem_data2[43]), .C2(n3242), .A(n1686), .B(n1687), .ZN(
        n1670) );
  AOI211_X2 U477 ( .C1(n3272), .C2(n1672), .A(n1673), .B(n1674), .ZN(n1671) );
  AOI211_X2 U480 ( .C1(ymem_data2[42]), .C2(n3242), .A(n1667), .B(n1668), .ZN(
        n1651) );
  AOI211_X2 U481 ( .C1(n3272), .C2(n1653), .A(n1654), .B(n1655), .ZN(n1652) );
  AOI211_X2 U484 ( .C1(ymem_data2[41]), .C2(n866), .A(n1648), .B(n1649), .ZN(
        n1632) );
  AOI211_X2 U486 ( .C1(n3272), .C2(n1634), .A(n1635), .B(n1636), .ZN(n1633) );
  AOI211_X2 U487 ( .C1(ymem_data2[40]), .C2(n866), .A(n1629), .B(n1630), .ZN(
        n1613) );
  AOI211_X2 U492 ( .C1(n3272), .C2(n1615), .A(n1616), .B(n1617), .ZN(n1614) );
  AOI211_X2 U497 ( .C1(ymem_data2[39]), .C2(n866), .A(n1610), .B(n1611), .ZN(
        n1594) );
  AOI211_X2 U500 ( .C1(n3272), .C2(n1596), .A(n1597), .B(n1598), .ZN(n1595) );
  AOI211_X2 U501 ( .C1(ymem_data2[38]), .C2(n866), .A(n1591), .B(n1592), .ZN(
        n1575) );
  AOI211_X2 U504 ( .C1(n3272), .C2(n1577), .A(n1578), .B(n1579), .ZN(n1576) );
  AOI211_X2 U506 ( .C1(ymem_data2[37]), .C2(n866), .A(n1572), .B(n1573), .ZN(
        n1556) );
  AOI211_X2 U507 ( .C1(n3272), .C2(n1558), .A(n1559), .B(n1560), .ZN(n1557) );
  AOI211_X2 U512 ( .C1(ymem_data2[36]), .C2(n866), .A(n1553), .B(n1554), .ZN(
        n1537) );
  AOI211_X2 U517 ( .C1(n3272), .C2(n1539), .A(n1540), .B(n1541), .ZN(n1538) );
  AOI211_X2 U520 ( .C1(ymem_data2[47]), .C2(n866), .A(n1773), .B(n1774), .ZN(
        n1746) );
  AOI211_X2 U521 ( .C1(n3272), .C2(n1748), .A(n1749), .B(n1750), .ZN(n1747) );
  AOI21_X2 U524 ( .B1(n1732), .B2(n1733), .A(n3200), .ZN(n1731) );
  AOI21_X2 U526 ( .B1(n1713), .B2(n1714), .A(n3200), .ZN(n1712) );
  AOI21_X2 U527 ( .B1(n1694), .B2(n1695), .A(n3200), .ZN(n1693) );
  AOI21_X2 U532 ( .B1(n1675), .B2(n1676), .A(n3200), .ZN(n1674) );
  AOI21_X2 U537 ( .B1(n1656), .B2(n1657), .A(n3200), .ZN(n1655) );
  AOI21_X2 U540 ( .B1(n1637), .B2(n1638), .A(n3200), .ZN(n1636) );
  AOI21_X2 U541 ( .B1(n1618), .B2(n1619), .A(n3200), .ZN(n1617) );
  AOI21_X2 U544 ( .B1(n1599), .B2(n1600), .A(n3200), .ZN(n1598) );
  AOI21_X2 U546 ( .B1(n1580), .B2(n1581), .A(n3200), .ZN(n1579) );
  AOI21_X2 U547 ( .B1(n1561), .B2(n1562), .A(n3200), .ZN(n1560) );
  AOI21_X2 U552 ( .B1(n1542), .B2(n1543), .A(n3200), .ZN(n1541) );
  AOI21_X2 U557 ( .B1(n1523), .B2(n1524), .A(n3200), .ZN(n1522) );
  AOI21_X2 U560 ( .B1(n1751), .B2(n1752), .A(n3200), .ZN(n1750) );
  OAI222_X2 U561 ( .A1(n562), .A2(n3230), .B1(n626), .B2(n1810), .C1(n498), 
        .C2(n3227), .ZN(n2144) );
  OAI222_X2 U564 ( .A1(n561), .A2(n3230), .B1(n625), .B2(n1810), .C1(n497), 
        .C2(n3227), .ZN(n2136) );
  OAI222_X2 U566 ( .A1(n560), .A2(n3231), .B1(n624), .B2(n3228), .C1(n496), 
        .C2(n3227), .ZN(n2059) );
  OAI222_X2 U567 ( .A1(n559), .A2(n3231), .B1(n623), .B2(n3228), .C1(n495), 
        .C2(n3227), .ZN(n1982) );
  OAI222_X2 U572 ( .A1(n558), .A2(n3231), .B1(n622), .B2(n1810), .C1(n494), 
        .C2(n3227), .ZN(n1905) );
  OAI222_X2 U577 ( .A1(n557), .A2(n3230), .B1(n621), .B2(n3228), .C1(n493), 
        .C2(n3227), .ZN(n1842) );
  OAI222_X2 U580 ( .A1(n556), .A2(n3230), .B1(n620), .B2(n3228), .C1(n492), 
        .C2(n3227), .ZN(n1835) );
  OAI222_X2 U581 ( .A1(n555), .A2(n3231), .B1(n619), .B2(n1810), .C1(n491), 
        .C2(n1811), .ZN(n1828) );
  OAI222_X2 U587 ( .A1(n552), .A2(n3230), .B1(n616), .B2(n1810), .C1(n488), 
        .C2(n3227), .ZN(n2129) );
  OAI222_X2 U592 ( .A1(n551), .A2(n3230), .B1(n615), .B2(n1810), .C1(n487), 
        .C2(n3227), .ZN(n2122) );
  OAI222_X2 U597 ( .A1(n550), .A2(n3230), .B1(n614), .B2(n1810), .C1(n486), 
        .C2(n3227), .ZN(n2115) );
  OAI222_X2 U600 ( .A1(n549), .A2(n3230), .B1(n613), .B2(n1810), .C1(n485), 
        .C2(n3227), .ZN(n2108) );
  OAI222_X2 U601 ( .A1(n548), .A2(n3230), .B1(n612), .B2(n3228), .C1(n484), 
        .C2(n1811), .ZN(n2101) );
  OAI222_X2 U604 ( .A1(n547), .A2(n3230), .B1(n611), .B2(n3228), .C1(n483), 
        .C2(n1811), .ZN(n2094) );
  OAI222_X2 U607 ( .A1(n545), .A2(n3230), .B1(n609), .B2(n1810), .C1(n481), 
        .C2(n1811), .ZN(n2080) );
  OAI222_X2 U617 ( .A1(n543), .A2(n3230), .B1(n607), .B2(n1810), .C1(n479), 
        .C2(n1811), .ZN(n2066) );
  OAI222_X2 U620 ( .A1(n542), .A2(n3231), .B1(n606), .B2(n3228), .C1(n478), 
        .C2(n3227), .ZN(n2052) );
  OAI222_X2 U621 ( .A1(n541), .A2(n3231), .B1(n605), .B2(n3228), .C1(n477), 
        .C2(n3227), .ZN(n2045) );
  OAI222_X2 U624 ( .A1(n540), .A2(n3231), .B1(n604), .B2(n3228), .C1(n476), 
        .C2(n3227), .ZN(n2038) );
  OAI222_X2 U626 ( .A1(n539), .A2(n3231), .B1(n603), .B2(n3228), .C1(n475), 
        .C2(n3227), .ZN(n2031) );
  OAI222_X2 U627 ( .A1(n538), .A2(n3231), .B1(n602), .B2(n3228), .C1(n474), 
        .C2(n3227), .ZN(n2024) );
  OAI222_X2 U632 ( .A1(n537), .A2(n3231), .B1(n601), .B2(n3228), .C1(n473), 
        .C2(n3227), .ZN(n2017) );
  OAI222_X2 U637 ( .A1(n536), .A2(n3231), .B1(n600), .B2(n3228), .C1(n472), 
        .C2(n3227), .ZN(n2010) );
  OAI222_X2 U640 ( .A1(n535), .A2(n3231), .B1(n599), .B2(n3228), .C1(n471), 
        .C2(n3227), .ZN(n2003) );
  OAI222_X2 U641 ( .A1(n534), .A2(n3231), .B1(n598), .B2(n3228), .C1(n470), 
        .C2(n3227), .ZN(n1996) );
  OAI222_X2 U644 ( .A1(n533), .A2(n3231), .B1(n597), .B2(n3228), .C1(n469), 
        .C2(n3227), .ZN(n1989) );
  OAI222_X2 U647 ( .A1(n531), .A2(n3230), .B1(n595), .B2(n3228), .C1(n467), 
        .C2(n1811), .ZN(n1968) );
  OAI222_X2 U652 ( .A1(n530), .A2(n3231), .B1(n594), .B2(n3228), .C1(n466), 
        .C2(n1811), .ZN(n1961) );
  OAI222_X2 U657 ( .A1(n529), .A2(n3230), .B1(n593), .B2(n3228), .C1(n465), 
        .C2(n1811), .ZN(n1954) );
  OAI222_X2 U660 ( .A1(n528), .A2(n3231), .B1(n592), .B2(n3228), .C1(n464), 
        .C2(n1811), .ZN(n1947) );
  OAI222_X2 U661 ( .A1(n527), .A2(n3230), .B1(n591), .B2(n3228), .C1(n463), 
        .C2(n1811), .ZN(n1940) );
  OAI222_X2 U664 ( .A1(n526), .A2(n3231), .B1(n590), .B2(n3228), .C1(n462), 
        .C2(n1811), .ZN(n1933) );
  OAI222_X2 U666 ( .A1(n525), .A2(n3230), .B1(n589), .B2(n3228), .C1(n461), 
        .C2(n1811), .ZN(n1926) );
  OAI222_X2 U667 ( .A1(n524), .A2(n3231), .B1(n588), .B2(n3228), .C1(n460), 
        .C2(n1811), .ZN(n1919) );
  OAI222_X2 U672 ( .A1(n523), .A2(n3230), .B1(n587), .B2(n3228), .C1(n459), 
        .C2(n1811), .ZN(n1912) );
  OAI222_X2 U677 ( .A1(n522), .A2(n3231), .B1(n586), .B2(n3228), .C1(n458), 
        .C2(n1811), .ZN(n1898) );
  OAI222_X2 U680 ( .A1(n521), .A2(n3231), .B1(n585), .B2(n1810), .C1(n457), 
        .C2(n1811), .ZN(n1891) );
  OAI222_X2 U681 ( .A1(n520), .A2(n3231), .B1(n584), .B2(n1810), .C1(n456), 
        .C2(n1811), .ZN(n1884) );
  OAI222_X2 U684 ( .A1(n519), .A2(n3230), .B1(n583), .B2(n1810), .C1(n455), 
        .C2(n3227), .ZN(n1877) );
  OAI222_X2 U686 ( .A1(n518), .A2(n3230), .B1(n582), .B2(n1810), .C1(n454), 
        .C2(n3227), .ZN(n1870) );
  OAI222_X2 U687 ( .A1(n517), .A2(n3231), .B1(n581), .B2(n1810), .C1(n453), 
        .C2(n3227), .ZN(n1863) );
  OAI222_X2 U692 ( .A1(n516), .A2(n3230), .B1(n580), .B2(n1810), .C1(n452), 
        .C2(n3227), .ZN(n1856) );
  OAI222_X2 U697 ( .A1(n515), .A2(n3231), .B1(n579), .B2(n1810), .C1(n451), 
        .C2(n3227), .ZN(n1849) );
  OAI21_X2 U700 ( .B1(n2551), .B2(n2552), .A(n131), .ZN(n2550) );
  OAI21_X2 U701 ( .B1(n785), .B2(n786), .A(n787), .ZN(n2628) );
  OAI222_X2 U704 ( .A1(n3278), .A2(n748), .B1(n744), .B2(n795), .C1(n796), 
        .C2(n797), .ZN(n789) );
  AOI211_X2 U706 ( .C1(n3273), .C2(n1520), .A(n1521), .B(n1522), .ZN(n1519) );
  AOI211_X2 U707 ( .C1(ymem_data2[35]), .C2(n3242), .A(n1534), .B(n1535), .ZN(
        n1518) );
  AOI21_X2 U712 ( .B1(n1527), .B2(n1528), .A(n3201), .ZN(n1521) );
  AOI211_X2 U717 ( .C1(n3273), .C2(n1501), .A(n1502), .B(n1503), .ZN(n1500) );
  AOI211_X2 U720 ( .C1(ymem_data2[34]), .C2(n3242), .A(n1515), .B(n1516), .ZN(
        n1499) );
  AOI21_X2 U721 ( .B1(n1508), .B2(n1509), .A(n3201), .ZN(n1502) );
  AOI211_X2 U724 ( .C1(n3273), .C2(n1482), .A(n1483), .B(n1484), .ZN(n1481) );
  AOI211_X2 U726 ( .C1(ymem_data2[33]), .C2(n3242), .A(n1496), .B(n1497), .ZN(
        n1480) );
  AOI21_X2 U727 ( .B1(n1489), .B2(n1490), .A(n3201), .ZN(n1483) );
  AOI211_X2 U732 ( .C1(n3273), .C2(n1463), .A(n1464), .B(n1465), .ZN(n1462) );
  AOI211_X2 U737 ( .C1(ymem_data2[32]), .C2(n3242), .A(n1477), .B(n1478), .ZN(
        n1461) );
  AOI21_X2 U740 ( .B1(n1470), .B2(n1471), .A(n3201), .ZN(n1464) );
  AOI211_X2 U741 ( .C1(n3273), .C2(n1444), .A(n1445), .B(n1446), .ZN(n1443) );
  AOI211_X2 U744 ( .C1(ymem_data2[31]), .C2(n3242), .A(n1458), .B(n1459), .ZN(
        n1442) );
  AOI21_X2 U746 ( .B1(n1451), .B2(n1452), .A(n3201), .ZN(n1445) );
  AOI211_X2 U747 ( .C1(n3273), .C2(n1425), .A(n1426), .B(n1427), .ZN(n1424) );
  AOI211_X2 U752 ( .C1(ymem_data2[30]), .C2(n3242), .A(n1439), .B(n1440), .ZN(
        n1423) );
  AOI21_X2 U757 ( .B1(n1432), .B2(n1433), .A(n3201), .ZN(n1426) );
  AOI211_X2 U760 ( .C1(n3273), .C2(n1406), .A(n1407), .B(n1408), .ZN(n1405) );
  AOI211_X2 U761 ( .C1(ymem_data2[29]), .C2(n3242), .A(n1420), .B(n1421), .ZN(
        n1404) );
  AOI21_X2 U764 ( .B1(n1413), .B2(n1414), .A(n3201), .ZN(n1407) );
  AOI211_X2 U766 ( .C1(n3273), .C2(n1387), .A(n1388), .B(n1389), .ZN(n1386) );
  AOI211_X2 U767 ( .C1(ymem_data2[28]), .C2(n3242), .A(n1401), .B(n1402), .ZN(
        n1385) );
  AOI21_X2 U772 ( .B1(n1394), .B2(n1395), .A(n3201), .ZN(n1388) );
  AOI211_X2 U777 ( .C1(n3273), .C2(n1368), .A(n1369), .B(n1370), .ZN(n1367) );
  AOI211_X2 U780 ( .C1(ymem_data2[27]), .C2(n3242), .A(n1382), .B(n1383), .ZN(
        n1366) );
  AOI21_X2 U781 ( .B1(n1375), .B2(n1376), .A(n3201), .ZN(n1369) );
  AOI211_X2 U784 ( .C1(n3273), .C2(n1349), .A(n1350), .B(n1351), .ZN(n1348) );
  AOI211_X2 U786 ( .C1(ymem_data2[26]), .C2(n3242), .A(n1363), .B(n1364), .ZN(
        n1347) );
  AOI21_X2 U787 ( .B1(n1356), .B2(n1357), .A(n3201), .ZN(n1350) );
  AOI211_X2 U792 ( .C1(n3273), .C2(n1330), .A(n1331), .B(n1332), .ZN(n1329) );
  AOI211_X2 U797 ( .C1(ymem_data2[25]), .C2(n3242), .A(n1344), .B(n1345), .ZN(
        n1328) );
  AOI21_X2 U800 ( .B1(n1337), .B2(n1338), .A(n3201), .ZN(n1331) );
  AOI211_X2 U801 ( .C1(n3273), .C2(n1311), .A(n1312), .B(n1313), .ZN(n1310) );
  AOI211_X2 U804 ( .C1(ymem_data2[24]), .C2(n3242), .A(n1325), .B(n1326), .ZN(
        n1309) );
  AOI21_X2 U806 ( .B1(n1318), .B2(n1319), .A(n3201), .ZN(n1312) );
  AOI211_X2 U807 ( .C1(n3273), .C2(n1292), .A(n1293), .B(n1294), .ZN(n1291) );
  AOI211_X2 U812 ( .C1(ymem_data2[23]), .C2(n3242), .A(n1306), .B(n1307), .ZN(
        n1290) );
  AOI21_X2 U817 ( .B1(n1299), .B2(n1300), .A(n3201), .ZN(n1293) );
  AOI211_X2 U820 ( .C1(n3272), .C2(n1273), .A(n1274), .B(n1275), .ZN(n1272) );
  AOI211_X2 U821 ( .C1(ymem_data2[22]), .C2(n866), .A(n1287), .B(n1288), .ZN(
        n1271) );
  AOI21_X2 U824 ( .B1(n1280), .B2(n1281), .A(n3201), .ZN(n1274) );
  AOI211_X2 U826 ( .C1(n3273), .C2(n1254), .A(n1255), .B(n1256), .ZN(n1253) );
  AOI211_X2 U827 ( .C1(ymem_data2[21]), .C2(n866), .A(n1268), .B(n1269), .ZN(
        n1252) );
  AOI21_X2 U832 ( .B1(n1261), .B2(n1262), .A(n3201), .ZN(n1255) );
  AOI211_X2 U837 ( .C1(n3272), .C2(n1235), .A(n1236), .B(n1237), .ZN(n1234) );
  AOI211_X2 U840 ( .C1(ymem_data2[20]), .C2(n3242), .A(n1249), .B(n1250), .ZN(
        n1233) );
  AOI21_X2 U841 ( .B1(n1242), .B2(n1243), .A(n3201), .ZN(n1236) );
  AOI211_X2 U844 ( .C1(n3273), .C2(n1216), .A(n1217), .B(n1218), .ZN(n1215) );
  AOI211_X2 U846 ( .C1(ymem_data2[19]), .C2(n3242), .A(n1230), .B(n1231), .ZN(
        n1214) );
  AOI21_X2 U847 ( .B1(n1223), .B2(n1224), .A(n3201), .ZN(n1217) );
  AOI211_X2 U852 ( .C1(n3272), .C2(n1197), .A(n1198), .B(n1199), .ZN(n1196) );
  AOI211_X2 U857 ( .C1(ymem_data2[18]), .C2(n3242), .A(n1211), .B(n1212), .ZN(
        n1195) );
  AOI21_X2 U860 ( .B1(n1204), .B2(n1205), .A(n3201), .ZN(n1198) );
  AOI211_X2 U861 ( .C1(n3273), .C2(n1178), .A(n1179), .B(n1180), .ZN(n1177) );
  AOI211_X2 U864 ( .C1(ymem_data2[17]), .C2(n3242), .A(n1192), .B(n1193), .ZN(
        n1176) );
  AOI21_X2 U866 ( .B1(n1185), .B2(n1186), .A(n3201), .ZN(n1179) );
  AOI211_X2 U867 ( .C1(n3272), .C2(n1159), .A(n1160), .B(n1161), .ZN(n1158) );
  AOI211_X2 U872 ( .C1(ymem_data2[16]), .C2(n3242), .A(n1173), .B(n1174), .ZN(
        n1157) );
  AOI21_X2 U877 ( .B1(n1166), .B2(n1167), .A(n3201), .ZN(n1160) );
  AOI211_X2 U880 ( .C1(n3273), .C2(n1140), .A(n1141), .B(n1142), .ZN(n1139) );
  AOI211_X2 U881 ( .C1(ymem_data2[15]), .C2(n3242), .A(n1154), .B(n1155), .ZN(
        n1138) );
  AOI21_X2 U884 ( .B1(n1147), .B2(n1148), .A(n3201), .ZN(n1141) );
  AOI211_X2 U886 ( .C1(n3272), .C2(n1121), .A(n1122), .B(n1123), .ZN(n1120) );
  AOI211_X2 U887 ( .C1(ymem_data2[14]), .C2(n3242), .A(n1135), .B(n1136), .ZN(
        n1119) );
  AOI21_X2 U892 ( .B1(n1128), .B2(n1129), .A(n3201), .ZN(n1122) );
  AOI211_X2 U897 ( .C1(n3273), .C2(n1102), .A(n1103), .B(n1104), .ZN(n1101) );
  AOI211_X2 U900 ( .C1(ymem_data2[13]), .C2(n3242), .A(n1116), .B(n1117), .ZN(
        n1100) );
  AOI21_X2 U901 ( .B1(n1109), .B2(n1110), .A(n3201), .ZN(n1103) );
  AOI211_X2 U904 ( .C1(n3273), .C2(n1083), .A(n1084), .B(n1085), .ZN(n1082) );
  AOI211_X2 U906 ( .C1(ymem_data2[12]), .C2(n3242), .A(n1097), .B(n1098), .ZN(
        n1081) );
  AOI21_X2 U907 ( .B1(n1090), .B2(n1091), .A(n3201), .ZN(n1084) );
  AOI211_X2 U912 ( .C1(n3273), .C2(n1064), .A(n1065), .B(n1066), .ZN(n1063) );
  AOI211_X2 U917 ( .C1(ymem_data2[11]), .C2(n866), .A(n1078), .B(n1079), .ZN(
        n1062) );
  AOI21_X2 U920 ( .B1(n1071), .B2(n1072), .A(n3201), .ZN(n1065) );
  AOI211_X2 U921 ( .C1(n3272), .C2(n1045), .A(n1046), .B(n1047), .ZN(n1044) );
  AOI211_X2 U924 ( .C1(ymem_data2[10]), .C2(n866), .A(n1059), .B(n1060), .ZN(
        n1043) );
  AOI21_X2 U926 ( .B1(n1052), .B2(n1053), .A(n3201), .ZN(n1046) );
  AOI211_X2 U927 ( .C1(n3272), .C2(n1026), .A(n1027), .B(n1028), .ZN(n1025) );
  AOI211_X2 U932 ( .C1(ymem_data2[9]), .C2(n866), .A(n1040), .B(n1041), .ZN(
        n1024) );
  AOI21_X2 U937 ( .B1(n1033), .B2(n1034), .A(n3201), .ZN(n1027) );
  AOI211_X2 U940 ( .C1(n3273), .C2(n1007), .A(n1008), .B(n1009), .ZN(n1006) );
  AOI211_X2 U941 ( .C1(ymem_data2[8]), .C2(n3242), .A(n1021), .B(n1022), .ZN(
        n1005) );
  AOI21_X2 U944 ( .B1(n1014), .B2(n1015), .A(n3201), .ZN(n1008) );
  AOI211_X2 U946 ( .C1(n3272), .C2(n988), .A(n989), .B(n990), .ZN(n987) );
  AOI211_X2 U947 ( .C1(ymem_data2[7]), .C2(n3242), .A(n1002), .B(n1003), .ZN(
        n986) );
  AOI21_X2 U952 ( .B1(n995), .B2(n996), .A(n3201), .ZN(n989) );
  AOI211_X2 U957 ( .C1(n3272), .C2(n969), .A(n970), .B(n971), .ZN(n968) );
  AOI211_X2 U960 ( .C1(ymem_data2[6]), .C2(n3242), .A(n983), .B(n984), .ZN(
        n967) );
  AOI21_X2 U961 ( .B1(n976), .B2(n977), .A(n3201), .ZN(n970) );
  AOI211_X2 U964 ( .C1(n3273), .C2(n950), .A(n951), .B(n952), .ZN(n949) );
  AOI211_X2 U966 ( .C1(ymem_data2[5]), .C2(n3242), .A(n964), .B(n965), .ZN(
        n948) );
  AOI21_X2 U967 ( .B1(n957), .B2(n958), .A(n3201), .ZN(n951) );
  AOI211_X2 U972 ( .C1(n3273), .C2(n931), .A(n932), .B(n933), .ZN(n930) );
  AOI211_X2 U977 ( .C1(ymem_data2[4]), .C2(n866), .A(n945), .B(n946), .ZN(n929) );
  AOI21_X2 U980 ( .B1(n938), .B2(n939), .A(n3201), .ZN(n932) );
  AOI211_X2 U981 ( .C1(n3272), .C2(n912), .A(n913), .B(n914), .ZN(n911) );
  AOI211_X2 U984 ( .C1(ymem_data2[3]), .C2(n866), .A(n926), .B(n927), .ZN(n910) );
  AOI21_X2 U986 ( .B1(n919), .B2(n920), .A(n3201), .ZN(n913) );
  AOI211_X2 U987 ( .C1(n3273), .C2(n893), .A(n894), .B(n895), .ZN(n892) );
  AOI211_X2 U992 ( .C1(ymem_data2[2]), .C2(n866), .A(n907), .B(n908), .ZN(n891) );
  AOI21_X2 U997 ( .B1(n900), .B2(n901), .A(n3201), .ZN(n894) );
  AOI211_X2 U1000 ( .C1(n3272), .C2(n874), .A(n875), .B(n876), .ZN(n873) );
  AOI211_X2 U1001 ( .C1(ymem_data2[1]), .C2(n866), .A(n888), .B(n889), .ZN(
        n872) );
  AOI21_X2 U1004 ( .B1(n881), .B2(n882), .A(n3201), .ZN(n875) );
  AOI211_X2 U1006 ( .C1(n3272), .C2(n837), .A(n838), .B(n839), .ZN(n835) );
  AOI211_X2 U1007 ( .C1(ymem_data2[0]), .C2(n866), .A(n867), .B(n868), .ZN(
        n832) );
  AOI21_X2 U1012 ( .B1(n845), .B2(n846), .A(n3201), .ZN(n838) );
  OAI211_X2 U1017 ( .C1(ymem_data1[255]), .C2(n129), .A(n2521), .B(n2522), 
        .ZN(n2512) );
  OAI211_X2 U1020 ( .C1(n3299), .C2(n580), .A(n1740), .B(n1741), .ZN(n1729) );
  AOI22_X2 U1021 ( .A1(ymem_data2[174]), .A2(n3246), .B1(ymem_data2[110]), 
        .B2(n865), .ZN(n1740) );
  OAI211_X2 U1024 ( .C1(n3299), .C2(n581), .A(n1721), .B(n1722), .ZN(n1710) );
  AOI22_X2 U1026 ( .A1(ymem_data2[173]), .A2(n3246), .B1(ymem_data2[109]), 
        .B2(n865), .ZN(n1721) );
  OAI211_X2 U1027 ( .C1(n3299), .C2(n582), .A(n1702), .B(n1703), .ZN(n1691) );
  AOI22_X2 U1032 ( .A1(ymem_data2[172]), .A2(n3246), .B1(ymem_data2[108]), 
        .B2(n3244), .ZN(n1702) );
  OAI211_X2 U1037 ( .C1(n3299), .C2(n583), .A(n1683), .B(n1684), .ZN(n1672) );
  AOI22_X2 U1040 ( .A1(ymem_data2[171]), .A2(n3246), .B1(ymem_data2[107]), 
        .B2(n3244), .ZN(n1683) );
  OAI211_X2 U1041 ( .C1(n3299), .C2(n584), .A(n1664), .B(n1665), .ZN(n1653) );
  AOI22_X2 U1044 ( .A1(ymem_data2[170]), .A2(n3246), .B1(ymem_data2[106]), 
        .B2(n865), .ZN(n1664) );
  OAI211_X2 U1046 ( .C1(n3299), .C2(n585), .A(n1645), .B(n1646), .ZN(n1634) );
  AOI22_X2 U1047 ( .A1(ymem_data2[169]), .A2(n3246), .B1(ymem_data2[105]), 
        .B2(n865), .ZN(n1645) );
  OAI211_X2 U1052 ( .C1(n3299), .C2(n586), .A(n1626), .B(n1627), .ZN(n1615) );
  AOI22_X2 U1057 ( .A1(ymem_data2[168]), .A2(n3246), .B1(ymem_data2[104]), 
        .B2(n865), .ZN(n1626) );
  OAI211_X2 U1060 ( .C1(n3299), .C2(n587), .A(n1607), .B(n1608), .ZN(n1596) );
  AOI22_X2 U1061 ( .A1(ymem_data2[167]), .A2(n3246), .B1(ymem_data2[103]), 
        .B2(n865), .ZN(n1607) );
  OAI211_X2 U1064 ( .C1(n3299), .C2(n588), .A(n1588), .B(n1589), .ZN(n1577) );
  AOI22_X2 U1066 ( .A1(ymem_data2[166]), .A2(n3246), .B1(ymem_data2[102]), 
        .B2(n865), .ZN(n1588) );
  OAI211_X2 U1067 ( .C1(n3299), .C2(n589), .A(n1569), .B(n1570), .ZN(n1558) );
  AOI22_X2 U1072 ( .A1(ymem_data2[165]), .A2(n3246), .B1(ymem_data2[101]), 
        .B2(n3244), .ZN(n1569) );
  OAI211_X2 U1077 ( .C1(n3299), .C2(n590), .A(n1550), .B(n1551), .ZN(n1539) );
  AOI22_X2 U1080 ( .A1(ymem_data2[164]), .A2(n3246), .B1(ymem_data2[100]), 
        .B2(n865), .ZN(n1550) );
  OAI211_X2 U1081 ( .C1(n3299), .C2(n579), .A(n1760), .B(n1761), .ZN(n1748) );
  AOI22_X2 U1084 ( .A1(ymem_data2[175]), .A2(n3246), .B1(ymem_data2[111]), 
        .B2(n865), .ZN(n1760) );
  AOI22_X2 U1086 ( .A1(ymem_data2[50]), .A2(n2472), .B1(ymem_data1[178]), .B2(
        n3287), .ZN(n2474) );
  AOI22_X2 U1087 ( .A1(ymem_data2[49]), .A2(n2472), .B1(ymem_data1[177]), .B2(
        n3287), .ZN(n2475) );
  AOI22_X2 U1088 ( .A1(ymem_data2[48]), .A2(n2472), .B1(ymem_data1[176]), .B2(
        n3287), .ZN(n2476) );
  AOI22_X2 U1091 ( .A1(ymem_data2[51]), .A2(n2472), .B1(ymem_data1[179]), .B2(
        n3287), .ZN(n2471) );
  AOI22_X2 U1092 ( .A1(ymem_data2[55]), .A2(n2472), .B1(ymem_data1[183]), .B2(
        n3287), .ZN(n2481) );
  AOI22_X2 U1094 ( .A1(ymem_data2[54]), .A2(n2472), .B1(ymem_data1[182]), .B2(
        n3287), .ZN(n2482) );
  AOI22_X2 U1098 ( .A1(ymem_data2[63]), .A2(n2472), .B1(ymem_data1[191]), .B2(
        n3287), .ZN(n2497) );
  AOI222_X1 U1100 ( .A1(ymem_data1[112]), .A2(n150), .B1(ymem_data1[240]), 
        .B2(n765), .C1(ymem_data1[48]), .C2(n3291), .ZN(n2524) );
  AOI22_X2 U1101 ( .A1(ymem_data1[252]), .A2(n125), .B1(ymem_data1[253]), .B2(
        n124), .ZN(n2560) );
  AOI222_X1 U1106 ( .A1(ymem_data1[115]), .A2(n150), .B1(ymem_data1[243]), 
        .B2(n765), .C1(ymem_data1[51]), .C2(n3291), .ZN(n2516) );
  OAI211_X2 U1109 ( .C1(n3299), .C2(n591), .A(n1531), .B(n1532), .ZN(n1520) );
  AOI22_X2 U1111 ( .A1(ymem_data2[163]), .A2(n3246), .B1(ymem_data2[99]), .B2(
        n3244), .ZN(n1531) );
  OAI211_X2 U1113 ( .C1(n3299), .C2(n592), .A(n1512), .B(n1513), .ZN(n1501) );
  AOI22_X2 U1114 ( .A1(ymem_data2[162]), .A2(n3246), .B1(ymem_data2[98]), .B2(
        n3244), .ZN(n1512) );
  OAI211_X2 U1116 ( .C1(n3299), .C2(n593), .A(n1493), .B(n1494), .ZN(n1482) );
  AOI22_X2 U1121 ( .A1(ymem_data2[161]), .A2(n3246), .B1(ymem_data2[97]), .B2(
        n3244), .ZN(n1493) );
  OAI211_X2 U1123 ( .C1(n3299), .C2(n594), .A(n1474), .B(n1475), .ZN(n1463) );
  AOI22_X2 U1124 ( .A1(ymem_data2[160]), .A2(n3246), .B1(ymem_data2[96]), .B2(
        n3244), .ZN(n1474) );
  OAI211_X2 U1126 ( .C1(n3299), .C2(n601), .A(n1341), .B(n1342), .ZN(n1330) );
  AOI22_X2 U1129 ( .A1(ymem_data2[153]), .A2(n3246), .B1(ymem_data2[89]), .B2(
        n3244), .ZN(n1341) );
  OAI211_X2 U1140 ( .C1(n3299), .C2(n602), .A(n1322), .B(n1323), .ZN(n1311) );
  AOI22_X2 U1146 ( .A1(ymem_data2[152]), .A2(n3246), .B1(ymem_data2[88]), .B2(
        n3244), .ZN(n1322) );
  OAI211_X2 U1148 ( .C1(n3299), .C2(n603), .A(n1303), .B(n1304), .ZN(n1292) );
  AOI22_X2 U1152 ( .A1(ymem_data2[151]), .A2(n864), .B1(ymem_data2[87]), .B2(
        n3244), .ZN(n1303) );
  OAI211_X2 U1159 ( .C1(n3299), .C2(n604), .A(n1284), .B(n1285), .ZN(n1273) );
  AOI22_X2 U1161 ( .A1(ymem_data2[150]), .A2(n864), .B1(ymem_data2[86]), .B2(
        n3244), .ZN(n1284) );
  OAI211_X2 U1162 ( .C1(n3299), .C2(n605), .A(n1265), .B(n1266), .ZN(n1254) );
  AOI22_X2 U1165 ( .A1(ymem_data2[149]), .A2(n864), .B1(ymem_data2[85]), .B2(
        n3244), .ZN(n1265) );
  OAI211_X2 U1167 ( .C1(n3299), .C2(n606), .A(n1246), .B(n1247), .ZN(n1235) );
  AOI22_X2 U1170 ( .A1(ymem_data2[148]), .A2(n864), .B1(ymem_data2[84]), .B2(
        n3244), .ZN(n1246) );
  OAI211_X2 U1172 ( .C1(n3299), .C2(n607), .A(n1227), .B(n1228), .ZN(n1216) );
  AOI22_X2 U1173 ( .A1(ymem_data2[147]), .A2(n864), .B1(ymem_data2[83]), .B2(
        n3244), .ZN(n1227) );
  OAI211_X2 U1175 ( .C1(n3299), .C2(n608), .A(n1208), .B(n1209), .ZN(n1197) );
  AOI22_X2 U1177 ( .A1(ymem_data2[146]), .A2(n864), .B1(ymem_data2[82]), .B2(
        n3244), .ZN(n1208) );
  OAI211_X2 U1180 ( .C1(n3299), .C2(n609), .A(n1189), .B(n1190), .ZN(n1178) );
  AOI22_X2 U1181 ( .A1(ymem_data2[145]), .A2(n864), .B1(ymem_data2[81]), .B2(
        n3244), .ZN(n1189) );
  OAI211_X2 U1183 ( .C1(n3299), .C2(n610), .A(n1170), .B(n1171), .ZN(n1159) );
  AOI22_X2 U1185 ( .A1(ymem_data2[144]), .A2(n864), .B1(ymem_data2[80]), .B2(
        n3244), .ZN(n1170) );
  OAI211_X2 U1188 ( .C1(n3299), .C2(n617), .A(n1037), .B(n1038), .ZN(n1026) );
  AOI22_X2 U1189 ( .A1(ymem_data2[137]), .A2(n3246), .B1(ymem_data2[73]), .B2(
        n865), .ZN(n1037) );
  OAI211_X2 U1191 ( .C1(n3299), .C2(n618), .A(n1018), .B(n1019), .ZN(n1007) );
  AOI22_X2 U1193 ( .A1(ymem_data2[136]), .A2(n3246), .B1(ymem_data2[72]), .B2(
        n865), .ZN(n1018) );
  OAI211_X2 U1196 ( .C1(n3299), .C2(n619), .A(n999), .B(n1000), .ZN(n988) );
  AOI22_X2 U1197 ( .A1(ymem_data2[135]), .A2(n3246), .B1(ymem_data2[71]), .B2(
        n865), .ZN(n999) );
  OAI211_X2 U1199 ( .C1(n3299), .C2(n620), .A(n980), .B(n981), .ZN(n969) );
  AOI22_X2 U1201 ( .A1(ymem_data2[134]), .A2(n864), .B1(ymem_data2[70]), .B2(
        n865), .ZN(n980) );
  OAI211_X2 U1204 ( .C1(n3299), .C2(n621), .A(n961), .B(n962), .ZN(n950) );
  AOI22_X2 U1205 ( .A1(ymem_data2[133]), .A2(n3246), .B1(ymem_data2[69]), .B2(
        n865), .ZN(n961) );
  OAI211_X2 U1207 ( .C1(n3299), .C2(n622), .A(n942), .B(n943), .ZN(n931) );
  AOI22_X2 U1209 ( .A1(ymem_data2[132]), .A2(n3246), .B1(ymem_data2[68]), .B2(
        n3244), .ZN(n942) );
  OAI211_X2 U1212 ( .C1(n3299), .C2(n623), .A(n923), .B(n924), .ZN(n912) );
  AOI22_X2 U1213 ( .A1(ymem_data2[131]), .A2(n864), .B1(ymem_data2[67]), .B2(
        n865), .ZN(n923) );
  OAI211_X2 U1215 ( .C1(n3299), .C2(n624), .A(n904), .B(n905), .ZN(n893) );
  AOI22_X2 U1217 ( .A1(ymem_data2[130]), .A2(n864), .B1(ymem_data2[66]), .B2(
        n3244), .ZN(n904) );
  OAI211_X2 U1220 ( .C1(n3299), .C2(n625), .A(n885), .B(n886), .ZN(n874) );
  AOI22_X2 U1221 ( .A1(ymem_data2[129]), .A2(n864), .B1(ymem_data2[65]), .B2(
        n3244), .ZN(n885) );
  OAI211_X2 U1223 ( .C1(n3299), .C2(n626), .A(n858), .B(n859), .ZN(n837) );
  AOI22_X2 U1225 ( .A1(ymem_data2[128]), .A2(n864), .B1(ymem_data2[64]), .B2(
        n865), .ZN(n858) );
  OAI211_X2 U1228 ( .C1(n3299), .C2(n595), .A(n1455), .B(n1456), .ZN(n1444) );
  AOI22_X2 U1229 ( .A1(ymem_data2[159]), .A2(n3246), .B1(ymem_data2[95]), .B2(
        n3244), .ZN(n1455) );
  OAI211_X2 U1231 ( .C1(n3299), .C2(n596), .A(n1436), .B(n1437), .ZN(n1425) );
  AOI22_X2 U1233 ( .A1(ymem_data2[158]), .A2(n3246), .B1(ymem_data2[94]), .B2(
        n3244), .ZN(n1436) );
  OAI211_X2 U1236 ( .C1(n3299), .C2(n597), .A(n1417), .B(n1418), .ZN(n1406) );
  AOI22_X2 U1237 ( .A1(ymem_data2[157]), .A2(n3246), .B1(ymem_data2[93]), .B2(
        n3244), .ZN(n1417) );
  OAI211_X2 U1239 ( .C1(n3299), .C2(n598), .A(n1398), .B(n1399), .ZN(n1387) );
  AOI22_X2 U1241 ( .A1(ymem_data2[156]), .A2(n864), .B1(ymem_data2[92]), .B2(
        n3244), .ZN(n1398) );
  OAI211_X2 U1244 ( .C1(n3299), .C2(n599), .A(n1379), .B(n1380), .ZN(n1368) );
  AOI22_X2 U1245 ( .A1(ymem_data2[155]), .A2(n864), .B1(ymem_data2[91]), .B2(
        n3244), .ZN(n1379) );
  OAI211_X2 U1247 ( .C1(n3299), .C2(n600), .A(n1360), .B(n1361), .ZN(n1349) );
  AOI22_X2 U1249 ( .A1(ymem_data2[154]), .A2(n864), .B1(ymem_data2[90]), .B2(
        n3244), .ZN(n1360) );
  OAI211_X2 U1252 ( .C1(n3299), .C2(n611), .A(n1151), .B(n1152), .ZN(n1140) );
  AOI22_X2 U1253 ( .A1(ymem_data2[143]), .A2(n864), .B1(ymem_data2[79]), .B2(
        n865), .ZN(n1151) );
  OAI211_X2 U1255 ( .C1(n3299), .C2(n612), .A(n1132), .B(n1133), .ZN(n1121) );
  AOI22_X2 U1257 ( .A1(ymem_data2[142]), .A2(n864), .B1(ymem_data2[78]), .B2(
        n865), .ZN(n1132) );
  OAI211_X2 U1260 ( .C1(n3299), .C2(n613), .A(n1113), .B(n1114), .ZN(n1102) );
  AOI22_X2 U1261 ( .A1(ymem_data2[141]), .A2(n864), .B1(ymem_data2[77]), .B2(
        n865), .ZN(n1113) );
  OAI211_X2 U1263 ( .C1(n3299), .C2(n614), .A(n1094), .B(n1095), .ZN(n1083) );
  AOI22_X2 U1265 ( .A1(ymem_data2[140]), .A2(n864), .B1(ymem_data2[76]), .B2(
        n865), .ZN(n1094) );
  OAI211_X2 U1268 ( .C1(n3299), .C2(n615), .A(n1075), .B(n1076), .ZN(n1064) );
  AOI22_X2 U1269 ( .A1(ymem_data2[139]), .A2(n3246), .B1(ymem_data2[75]), .B2(
        n3244), .ZN(n1075) );
  OAI211_X2 U1271 ( .C1(n3299), .C2(n616), .A(n1056), .B(n1057), .ZN(n1045) );
  AOI22_X2 U1273 ( .A1(ymem_data2[138]), .A2(n864), .B1(ymem_data2[74]), .B2(
        n3244), .ZN(n1056) );
  AOI222_X1 U1276 ( .A1(ymem_data1[119]), .A2(n150), .B1(ymem_data1[247]), 
        .B2(n765), .C1(ymem_data1[55]), .C2(n3291), .ZN(n2544) );
  AOI222_X1 U1277 ( .A1(ymem_data1[116]), .A2(n150), .B1(ymem_data1[244]), 
        .B2(n765), .C1(ymem_data1[52]), .C2(n3291), .ZN(n2535) );
  AOI21_X2 U1279 ( .B1(n1504), .B2(n1505), .A(n3200), .ZN(n1503) );
  AOI21_X2 U1281 ( .B1(n1485), .B2(n1486), .A(n3200), .ZN(n1484) );
  AOI21_X2 U1284 ( .B1(n1466), .B2(n1467), .A(n3200), .ZN(n1465) );
  AOI21_X2 U1285 ( .B1(n1447), .B2(n1448), .A(n3200), .ZN(n1446) );
  AOI21_X2 U1287 ( .B1(n1428), .B2(n1429), .A(n3200), .ZN(n1427) );
  AOI21_X2 U1289 ( .B1(n1409), .B2(n1410), .A(n3200), .ZN(n1408) );
  AOI21_X2 U1292 ( .B1(n1390), .B2(n1391), .A(n3200), .ZN(n1389) );
  AOI21_X2 U1293 ( .B1(n1371), .B2(n1372), .A(n3200), .ZN(n1370) );
  AOI21_X2 U1295 ( .B1(n1352), .B2(n1353), .A(n3200), .ZN(n1351) );
  AOI21_X2 U1297 ( .B1(n1333), .B2(n1334), .A(n3200), .ZN(n1332) );
  AOI21_X2 U1300 ( .B1(n1314), .B2(n1315), .A(n3200), .ZN(n1313) );
  AOI21_X2 U1301 ( .B1(n1295), .B2(n1296), .A(n3200), .ZN(n1294) );
  AOI21_X2 U1303 ( .B1(n1276), .B2(n1277), .A(n3200), .ZN(n1275) );
  AOI21_X2 U1305 ( .B1(n1257), .B2(n1258), .A(n3200), .ZN(n1256) );
  AOI21_X2 U1308 ( .B1(n1238), .B2(n1239), .A(n3200), .ZN(n1237) );
  AOI21_X2 U1309 ( .B1(n1219), .B2(n1220), .A(n3200), .ZN(n1218) );
  AOI21_X2 U1311 ( .B1(n1200), .B2(n1201), .A(n3200), .ZN(n1199) );
  AOI21_X2 U1313 ( .B1(n1181), .B2(n1182), .A(n3200), .ZN(n1180) );
  AOI21_X2 U1316 ( .B1(n1162), .B2(n1163), .A(n3200), .ZN(n1161) );
  AOI21_X2 U1317 ( .B1(n1143), .B2(n1144), .A(n3200), .ZN(n1142) );
  AOI21_X2 U1319 ( .B1(n1124), .B2(n1125), .A(n3200), .ZN(n1123) );
  AOI21_X2 U1321 ( .B1(n1105), .B2(n1106), .A(n3200), .ZN(n1104) );
  AOI21_X2 U1324 ( .B1(n1086), .B2(n1087), .A(n3200), .ZN(n1085) );
  AOI21_X2 U1325 ( .B1(n1067), .B2(n1068), .A(n3200), .ZN(n1066) );
  AOI21_X2 U1327 ( .B1(n1048), .B2(n1049), .A(n3200), .ZN(n1047) );
  AOI21_X2 U1329 ( .B1(n1029), .B2(n1030), .A(n3200), .ZN(n1028) );
  AOI21_X2 U1332 ( .B1(n1010), .B2(n1011), .A(n3200), .ZN(n1009) );
  AOI21_X2 U1333 ( .B1(n991), .B2(n992), .A(n3200), .ZN(n990) );
  AOI21_X2 U1335 ( .B1(n972), .B2(n973), .A(n3200), .ZN(n971) );
  AOI21_X2 U1337 ( .B1(n953), .B2(n954), .A(n3200), .ZN(n952) );
  AOI21_X2 U1340 ( .B1(n934), .B2(n935), .A(n3200), .ZN(n933) );
  AOI21_X2 U1341 ( .B1(n915), .B2(n916), .A(n3200), .ZN(n914) );
  AOI21_X2 U1343 ( .B1(n896), .B2(n897), .A(n3200), .ZN(n895) );
  AOI21_X2 U1345 ( .B1(n877), .B2(n878), .A(n3200), .ZN(n876) );
  AOI21_X2 U1348 ( .B1(n840), .B2(n841), .A(n3200), .ZN(n839) );
  AOI21_X2 U1349 ( .B1(n1736), .B2(n1737), .A(n3201), .ZN(n1730) );
  AOI21_X2 U1351 ( .B1(n1717), .B2(n1718), .A(n3201), .ZN(n1711) );
  AOI21_X2 U1353 ( .B1(n1698), .B2(n1699), .A(n3201), .ZN(n1692) );
  AOI21_X2 U1356 ( .B1(n1679), .B2(n1680), .A(n3201), .ZN(n1673) );
  AOI21_X2 U1357 ( .B1(n1660), .B2(n1661), .A(n3201), .ZN(n1654) );
  AOI21_X2 U1359 ( .B1(n1641), .B2(n1642), .A(n3201), .ZN(n1635) );
  AOI21_X2 U1361 ( .B1(n1622), .B2(n1623), .A(n3201), .ZN(n1616) );
  AOI21_X2 U1364 ( .B1(n1603), .B2(n1604), .A(n3201), .ZN(n1597) );
  AOI21_X2 U1365 ( .B1(n1584), .B2(n1585), .A(n3201), .ZN(n1578) );
  AOI21_X2 U1367 ( .B1(n1565), .B2(n1566), .A(n3201), .ZN(n1559) );
  AOI21_X2 U1369 ( .B1(n1546), .B2(n1547), .A(n3201), .ZN(n1540) );
  AOI21_X2 U1372 ( .B1(n1756), .B2(n1757), .A(n3201), .ZN(n1749) );
  OAI211_X2 U1373 ( .C1(n633), .C2(n634), .A(n635), .B(n636), .ZN(n2617) );
  AOI22_X2 U1375 ( .A1(yAddrIn1[0]), .A2(n642), .B1(yAddrIn2[0]), .B2(n643), 
        .ZN(n635) );
  OAI211_X2 U1377 ( .C1(n647), .C2(n634), .A(n648), .B(n649), .ZN(n2618) );
  AOI22_X2 U1380 ( .A1(yAddrIn1[1]), .A2(n642), .B1(yAddrIn2[1]), .B2(n643), 
        .ZN(n648) );
  OAI211_X2 U1381 ( .C1(n651), .C2(n634), .A(n652), .B(n653), .ZN(n2619) );
  AOI22_X2 U1383 ( .A1(yAddrIn1[2]), .A2(n642), .B1(yAddrIn2[2]), .B2(n643), 
        .ZN(n652) );
  OAI211_X2 U1385 ( .C1(n655), .C2(n634), .A(n656), .B(n657), .ZN(n2620) );
  AOI22_X2 U1388 ( .A1(yAddrIn1[3]), .A2(n642), .B1(yAddrIn2[3]), .B2(n643), 
        .ZN(n656) );
  OAI211_X2 U1389 ( .C1(n659), .C2(n634), .A(n660), .B(n661), .ZN(n2621) );
  AOI22_X2 U1391 ( .A1(yAddrIn1[4]), .A2(n642), .B1(yAddrIn2[4]), .B2(n643), 
        .ZN(n660) );
  OAI211_X2 U1393 ( .C1(n663), .C2(n634), .A(n664), .B(n665), .ZN(n2622) );
  AOI22_X2 U1396 ( .A1(yAddrIn1[5]), .A2(n642), .B1(yAddrIn2[5]), .B2(n643), 
        .ZN(n664) );
  OAI211_X2 U1397 ( .C1(n667), .C2(n634), .A(n668), .B(n669), .ZN(n2623) );
  AOI22_X2 U1399 ( .A1(yAddrIn1[6]), .A2(n642), .B1(yAddrIn2[6]), .B2(n643), 
        .ZN(n668) );
  OAI211_X2 U1401 ( .C1(n671), .C2(n634), .A(n672), .B(n673), .ZN(n2624) );
  AOI22_X2 U1404 ( .A1(yAddrIn1[7]), .A2(n642), .B1(yAddrIn2[7]), .B2(n643), 
        .ZN(n672) );
  OAI211_X2 U1405 ( .C1(n675), .C2(n3219), .A(n676), .B(n677), .ZN(n2625) );
  AOI22_X2 U1407 ( .A1(yAddrIn1[8]), .A2(n642), .B1(yAddrIn2[8]), .B2(n643), 
        .ZN(n676) );
  OAI211_X2 U1409 ( .C1(n679), .C2(n634), .A(n680), .B(n681), .ZN(n2626) );
  AOI22_X2 U1412 ( .A1(yAddrIn1[9]), .A2(n642), .B1(yAddrIn2[9]), .B2(n643), 
        .ZN(n680) );
  OAI211_X2 U1413 ( .C1(n683), .C2(n634), .A(n684), .B(n685), .ZN(n2627) );
  AOI22_X2 U1415 ( .A1(yAddrIn1[10]), .A2(n642), .B1(yAddrIn2[10]), .B2(n643), 
        .ZN(n684) );
  AOI21_X2 U1417 ( .B1(n2138), .B2(n2139), .A(n3301), .ZN(U94_Z_0) );
  AOI222_X1 U1420 ( .A1(ymem_data1[0]), .A2(n3289), .B1(n3202), .B2(
        U72_DATA1_0), .C1(ymem_data1[64]), .C2(n3288), .ZN(n2139) );
  AOI21_X2 U1421 ( .B1(n2142), .B2(n2143), .A(n3286), .ZN(n2141) );
  AOI21_X2 U1423 ( .B1(n2131), .B2(n2132), .A(n3301), .ZN(U94_Z_1) );
  AOI222_X1 U1425 ( .A1(ymem_data1[1]), .A2(n3289), .B1(n3202), .B2(
        U72_DATA1_1), .C1(ymem_data1[65]), .C2(n3288), .ZN(n2132) );
  AOI21_X2 U1428 ( .B1(n2134), .B2(n2135), .A(n3286), .ZN(n2133) );
  AOI21_X2 U1429 ( .B1(n2054), .B2(n2055), .A(n3301), .ZN(U94_Z_2) );
  AOI222_X1 U1431 ( .A1(ymem_data1[2]), .A2(n628), .B1(n3202), .B2(U72_DATA1_2), .C1(ymem_data1[66]), .C2(n3288), .ZN(n2055) );
  AOI21_X2 U1433 ( .B1(n2057), .B2(n2058), .A(n3286), .ZN(n2056) );
  AOI21_X2 U1436 ( .B1(n1977), .B2(n1978), .A(n3300), .ZN(U94_Z_3) );
  AOI222_X1 U1437 ( .A1(ymem_data1[3]), .A2(n628), .B1(n3202), .B2(U72_DATA1_3), .C1(ymem_data1[67]), .C2(n3288), .ZN(n1978) );
  AOI21_X2 U1439 ( .B1(n1980), .B2(n1981), .A(n715), .ZN(n1979) );
  AOI21_X2 U1441 ( .B1(n1900), .B2(n1901), .A(n3300), .ZN(U94_Z_4) );
  AOI222_X1 U1444 ( .A1(ymem_data1[4]), .A2(n628), .B1(n3202), .B2(U72_DATA1_4), .C1(ymem_data1[68]), .C2(n3288), .ZN(n1901) );
  AOI21_X2 U1445 ( .B1(n1903), .B2(n1904), .A(n3286), .ZN(n1902) );
  AOI21_X2 U1447 ( .B1(n2124), .B2(n2125), .A(n3301), .ZN(U94_Z_10) );
  AOI222_X1 U1449 ( .A1(ymem_data1[10]), .A2(n3289), .B1(n3202), .B2(
        U72_DATA1_10), .C1(ymem_data1[74]), .C2(n3288), .ZN(n2125) );
  AOI21_X2 U1452 ( .B1(n2127), .B2(n2128), .A(n3286), .ZN(n2126) );
  AOI21_X2 U1453 ( .B1(n2117), .B2(n2118), .A(n3301), .ZN(U94_Z_11) );
  AOI222_X1 U1455 ( .A1(ymem_data1[11]), .A2(n3289), .B1(n3202), .B2(
        U72_DATA1_11), .C1(ymem_data1[75]), .C2(n3288), .ZN(n2118) );
  AOI21_X2 U1457 ( .B1(n2120), .B2(n2121), .A(n3286), .ZN(n2119) );
  AOI21_X2 U1460 ( .B1(n1837), .B2(n1838), .A(n3300), .ZN(U94_Z_5) );
  AOI222_X1 U1461 ( .A1(ymem_data1[5]), .A2(n628), .B1(n3202), .B2(U72_DATA1_5), .C1(ymem_data1[69]), .C2(n3288), .ZN(n1838) );
  AOI21_X2 U1463 ( .B1(n1840), .B2(n1841), .A(n3286), .ZN(n1839) );
  AOI21_X2 U1465 ( .B1(n1830), .B2(n1831), .A(n3300), .ZN(U94_Z_6) );
  AOI222_X1 U1468 ( .A1(ymem_data1[6]), .A2(n3289), .B1(n3202), .B2(
        U72_DATA1_6), .C1(ymem_data1[70]), .C2(n3288), .ZN(n1831) );
  AOI21_X2 U1469 ( .B1(n1833), .B2(n1834), .A(n3286), .ZN(n1832) );
  AOI21_X2 U1471 ( .B1(n1823), .B2(n1824), .A(n3300), .ZN(U94_Z_7) );
  AOI222_X1 U1473 ( .A1(ymem_data1[7]), .A2(n628), .B1(n3202), .B2(U72_DATA1_7), .C1(ymem_data1[71]), .C2(n3288), .ZN(n1824) );
  AOI21_X2 U1476 ( .B1(n1826), .B2(n1827), .A(n3286), .ZN(n1825) );
  AOI21_X2 U1477 ( .B1(n1816), .B2(n1817), .A(n3300), .ZN(U94_Z_8) );
  AOI222_X1 U1479 ( .A1(ymem_data1[8]), .A2(n628), .B1(n3202), .B2(U72_DATA1_8), .C1(ymem_data1[72]), .C2(n3288), .ZN(n1817) );
  AOI21_X2 U1481 ( .B1(n1819), .B2(n1820), .A(n3286), .ZN(n1818) );
  AOI21_X2 U1484 ( .B1(n1801), .B2(n1802), .A(n3300), .ZN(U94_Z_9) );
  AOI222_X1 U1485 ( .A1(ymem_data1[9]), .A2(n3289), .B1(n3202), .B2(
        U72_DATA1_9), .C1(ymem_data1[73]), .C2(n3288), .ZN(n1802) );
  AOI21_X2 U1487 ( .B1(n1804), .B2(n1805), .A(n3286), .ZN(n1803) );
  AOI21_X2 U1489 ( .B1(n2110), .B2(n2111), .A(n3301), .ZN(U94_Z_12) );
  AOI222_X1 U1492 ( .A1(ymem_data1[12]), .A2(n3289), .B1(n3202), .B2(
        U72_DATA1_12), .C1(ymem_data1[76]), .C2(n3288), .ZN(n2111) );
  AOI21_X2 U1493 ( .B1(n2113), .B2(n2114), .A(n3286), .ZN(n2112) );
  AOI21_X2 U1495 ( .B1(n2103), .B2(n2104), .A(n3301), .ZN(U94_Z_13) );
  AOI222_X1 U1497 ( .A1(ymem_data1[13]), .A2(n3289), .B1(n3202), .B2(
        U72_DATA1_13), .C1(ymem_data1[77]), .C2(n3288), .ZN(n2104) );
  AOI21_X2 U1500 ( .B1(n2106), .B2(n2107), .A(n3286), .ZN(n2105) );
  AOI21_X2 U1501 ( .B1(n2096), .B2(n2097), .A(n3301), .ZN(U94_Z_14) );
  AOI222_X1 U1503 ( .A1(ymem_data1[14]), .A2(n3289), .B1(n3202), .B2(
        U72_DATA1_14), .C1(ymem_data1[78]), .C2(n3288), .ZN(n2097) );
  AOI21_X2 U1505 ( .B1(n2099), .B2(n2100), .A(n3286), .ZN(n2098) );
  AOI21_X2 U1508 ( .B1(n2089), .B2(n2090), .A(n3301), .ZN(U94_Z_15) );
  AOI222_X1 U1509 ( .A1(ymem_data1[15]), .A2(n3289), .B1(n3202), .B2(
        U72_DATA1_15), .C1(ymem_data1[79]), .C2(n3288), .ZN(n2090) );
  AOI21_X2 U1511 ( .B1(n2092), .B2(n2093), .A(n3286), .ZN(n2091) );
  AOI21_X2 U1513 ( .B1(n2082), .B2(n2083), .A(n3300), .ZN(U94_Z_16) );
  AOI222_X1 U1516 ( .A1(ymem_data1[16]), .A2(n3289), .B1(n3202), .B2(
        U72_DATA1_16), .C1(ymem_data1[80]), .C2(n3288), .ZN(n2083) );
  AOI21_X2 U1517 ( .B1(n2085), .B2(n2086), .A(n3286), .ZN(n2084) );
  AOI21_X2 U1519 ( .B1(n2075), .B2(n2076), .A(n3300), .ZN(U94_Z_17) );
  AOI222_X1 U1521 ( .A1(ymem_data1[17]), .A2(n3289), .B1(n3202), .B2(
        U72_DATA1_17), .C1(ymem_data1[81]), .C2(n3288), .ZN(n2076) );
  AOI21_X2 U1524 ( .B1(n2078), .B2(n2079), .A(n3286), .ZN(n2077) );
  AOI21_X2 U1525 ( .B1(n2068), .B2(n2069), .A(n3300), .ZN(U94_Z_18) );
  AOI222_X1 U1527 ( .A1(ymem_data1[18]), .A2(n3289), .B1(n3202), .B2(
        U72_DATA1_18), .C1(ymem_data1[82]), .C2(n3288), .ZN(n2069) );
  AOI21_X2 U1529 ( .B1(n2071), .B2(n2072), .A(n3286), .ZN(n2070) );
  AOI21_X2 U1532 ( .B1(n2061), .B2(n2062), .A(n3300), .ZN(U94_Z_19) );
  AOI222_X1 U1533 ( .A1(ymem_data1[19]), .A2(n3289), .B1(n3202), .B2(
        U72_DATA1_19), .C1(ymem_data1[83]), .C2(n3288), .ZN(n2062) );
  AOI21_X2 U1535 ( .B1(n2064), .B2(n2065), .A(n3286), .ZN(n2063) );
  AOI21_X2 U1537 ( .B1(n2047), .B2(n2048), .A(n3300), .ZN(U94_Z_20) );
  AOI222_X1 U1540 ( .A1(ymem_data1[20]), .A2(n628), .B1(n3202), .B2(
        U72_DATA1_20), .C1(ymem_data1[84]), .C2(n3288), .ZN(n2048) );
  AOI21_X2 U1541 ( .B1(n2050), .B2(n2051), .A(n3286), .ZN(n2049) );
  AOI21_X2 U1543 ( .B1(n2040), .B2(n2041), .A(n3300), .ZN(U94_Z_21) );
  AOI222_X1 U1545 ( .A1(ymem_data1[21]), .A2(n628), .B1(n3202), .B2(
        U72_DATA1_21), .C1(ymem_data1[85]), .C2(n3288), .ZN(n2041) );
  AOI21_X2 U1548 ( .B1(n2043), .B2(n2044), .A(n3286), .ZN(n2042) );
  AOI21_X2 U1549 ( .B1(n2033), .B2(n2034), .A(n3300), .ZN(U94_Z_22) );
  AOI222_X1 U1550 ( .A1(ymem_data1[22]), .A2(n628), .B1(n3202), .B2(
        U72_DATA1_22), .C1(ymem_data1[86]), .C2(n3288), .ZN(n2034) );
  AOI21_X2 U1551 ( .B1(n2036), .B2(n2037), .A(n3286), .ZN(n2035) );
  AOI21_X2 U1554 ( .B1(n2026), .B2(n2027), .A(n3300), .ZN(U94_Z_23) );
  AOI222_X1 U1556 ( .A1(ymem_data1[23]), .A2(n628), .B1(n3202), .B2(
        U72_DATA1_23), .C1(ymem_data1[87]), .C2(n3288), .ZN(n2027) );
  AOI21_X2 U1565 ( .B1(n2019), .B2(n2020), .A(n3300), .ZN(U94_Z_24) );
  AOI222_X1 U1570 ( .A1(ymem_data1[24]), .A2(n628), .B1(n3202), .B2(
        U72_DATA1_24), .C1(ymem_data1[88]), .C2(n3288), .ZN(n2020) );
  AOI21_X2 U1571 ( .B1(n2022), .B2(n2023), .A(n3286), .ZN(n2021) );
  AOI21_X2 U1580 ( .B1(n2012), .B2(n2013), .A(n3300), .ZN(U94_Z_25) );
  AOI222_X1 U1583 ( .A1(ymem_data1[25]), .A2(n628), .B1(n3202), .B2(
        U72_DATA1_25), .C1(ymem_data1[89]), .C2(n3288), .ZN(n2013) );
  AOI21_X2 U1606 ( .B1(n2005), .B2(n2006), .A(n3300), .ZN(U94_Z_26) );
  AOI222_X1 U1607 ( .A1(ymem_data1[26]), .A2(n628), .B1(n3202), .B2(
        U72_DATA1_26), .C1(ymem_data1[90]), .C2(n3288), .ZN(n2006) );
  AOI21_X2 U1611 ( .B1(n2008), .B2(n2009), .A(n3286), .ZN(n2007) );
  AOI21_X2 U1613 ( .B1(n1998), .B2(n1999), .A(n3301), .ZN(U94_Z_27) );
  AOI222_X1 U1614 ( .A1(ymem_data1[27]), .A2(n628), .B1(n3202), .B2(
        U72_DATA1_27), .C1(ymem_data1[91]), .C2(n3288), .ZN(n1999) );
  AOI21_X2 U1640 ( .B1(n1991), .B2(n1992), .A(n3300), .ZN(U94_Z_28) );
  AOI222_X1 U1682 ( .A1(ymem_data1[28]), .A2(n628), .B1(n3202), .B2(
        U72_DATA1_28), .C1(ymem_data1[92]), .C2(n3288), .ZN(n1992) );
  AOI21_X2 U1687 ( .B1(n1994), .B2(n1995), .A(n3286), .ZN(n1993) );
  AOI21_X2 U1688 ( .B1(n1984), .B2(n1985), .A(n3300), .ZN(U94_Z_29) );
  AOI222_X1 U1691 ( .A1(ymem_data1[29]), .A2(n628), .B1(n3202), .B2(
        U72_DATA1_29), .C1(ymem_data1[93]), .C2(n3288), .ZN(n1985) );
  AOI21_X2 U1695 ( .B1(n1970), .B2(n1971), .A(n3300), .ZN(U94_Z_30) );
  AOI222_X1 U1696 ( .A1(ymem_data1[30]), .A2(n3289), .B1(n3202), .B2(
        U72_DATA1_30), .C1(ymem_data1[94]), .C2(n3288), .ZN(n1971) );
  AOI21_X2 U1699 ( .B1(n1973), .B2(n1974), .A(n3286), .ZN(n1972) );
  AOI21_X2 U1700 ( .B1(n1963), .B2(n1964), .A(n3300), .ZN(U94_Z_31) );
  AOI222_X1 U1704 ( .A1(ymem_data1[31]), .A2(n3289), .B1(n3202), .B2(
        U72_DATA1_31), .C1(ymem_data1[95]), .C2(n3288), .ZN(n1964) );
  AOI21_X2 U1708 ( .B1(n1956), .B2(n1957), .A(n3300), .ZN(U94_Z_32) );
  AOI222_X1 U1709 ( .A1(ymem_data1[32]), .A2(n3289), .B1(n3202), .B2(
        U72_DATA1_32), .C1(ymem_data1[96]), .C2(n3288), .ZN(n1957) );
  AOI21_X2 U1712 ( .B1(n1959), .B2(n1960), .A(n3286), .ZN(n1958) );
  AOI21_X2 U1713 ( .B1(n1949), .B2(n1950), .A(n3300), .ZN(U94_Z_33) );
  AOI222_X1 U1716 ( .A1(ymem_data1[33]), .A2(n628), .B1(n3202), .B2(
        U72_DATA1_33), .C1(ymem_data1[97]), .C2(n3288), .ZN(n1950) );
  AOI21_X2 U1717 ( .B1(n1952), .B2(n1953), .A(n715), .ZN(n1951) );
  AOI21_X2 U1721 ( .B1(n1942), .B2(n1943), .A(n3300), .ZN(U94_Z_34) );
  AOI222_X1 U1722 ( .A1(ymem_data1[34]), .A2(n628), .B1(n3202), .B2(
        U72_DATA1_34), .C1(ymem_data1[98]), .C2(n3288), .ZN(n1943) );
  AOI21_X2 U1725 ( .B1(n1945), .B2(n1946), .A(n3286), .ZN(n1944) );
  AOI21_X2 U1726 ( .B1(n1935), .B2(n1936), .A(n3300), .ZN(U94_Z_35) );
  AOI222_X1 U1729 ( .A1(ymem_data1[35]), .A2(n628), .B1(n3202), .B2(
        U72_DATA1_35), .C1(ymem_data1[99]), .C2(n3288), .ZN(n1936) );
  AOI21_X2 U1730 ( .B1(n1938), .B2(n1939), .A(n3286), .ZN(n1937) );
  AOI21_X2 U1733 ( .B1(n1928), .B2(n1929), .A(n3300), .ZN(U94_Z_36) );
  AOI222_X1 U1734 ( .A1(ymem_data1[36]), .A2(n628), .B1(n3202), .B2(
        U72_DATA1_36), .C1(ymem_data1[100]), .C2(n3288), .ZN(n1929) );
  AOI21_X2 U1738 ( .B1(n1931), .B2(n1932), .A(n3286), .ZN(n1930) );
  AOI21_X2 U1739 ( .B1(n1921), .B2(n1922), .A(n3300), .ZN(U94_Z_37) );
  AOI222_X1 U1742 ( .A1(ymem_data1[37]), .A2(n3289), .B1(n3202), .B2(
        U72_DATA1_37), .C1(ymem_data1[101]), .C2(n3288), .ZN(n1922) );
  AOI21_X2 U1743 ( .B1(n1924), .B2(n1925), .A(n3286), .ZN(n1923) );
  AOI21_X2 U1746 ( .B1(n1914), .B2(n1915), .A(n3300), .ZN(U94_Z_38) );
  AOI222_X1 U1747 ( .A1(ymem_data1[38]), .A2(n628), .B1(n3202), .B2(
        U72_DATA1_38), .C1(ymem_data1[102]), .C2(n3288), .ZN(n1915) );
  AOI21_X2 U1750 ( .B1(n1917), .B2(n1918), .A(n3286), .ZN(n1916) );
  AOI21_X2 U1751 ( .B1(n1907), .B2(n1908), .A(n3300), .ZN(U94_Z_39) );
  AOI222_X1 U1752 ( .A1(ymem_data1[39]), .A2(n628), .B1(n3202), .B2(
        U72_DATA1_39), .C1(ymem_data1[103]), .C2(n3288), .ZN(n1908) );
  AOI21_X2 U1754 ( .B1(n1910), .B2(n1911), .A(n3286), .ZN(n1909) );
  AOI21_X2 U1760 ( .B1(n1893), .B2(n1894), .A(n3300), .ZN(U94_Z_40) );
  AOI222_X1 U1762 ( .A1(ymem_data1[40]), .A2(n628), .B1(n3202), .B2(
        U72_DATA1_40), .C1(ymem_data1[104]), .C2(n3288), .ZN(n1894) );
  AOI21_X2 U1764 ( .B1(n1896), .B2(n1897), .A(n3286), .ZN(n1895) );
  AOI21_X2 U1766 ( .B1(n1886), .B2(n1887), .A(n3300), .ZN(U94_Z_41) );
  AOI222_X1 U1769 ( .A1(ymem_data1[41]), .A2(n628), .B1(n3202), .B2(
        U72_DATA1_41), .C1(ymem_data1[105]), .C2(n3288), .ZN(n1887) );
  AOI21_X2 U1771 ( .B1(n1889), .B2(n1890), .A(n3286), .ZN(n1888) );
  AOI21_X2 U1773 ( .B1(n1879), .B2(n1880), .A(n3300), .ZN(U94_Z_42) );
  AOI222_X1 U1775 ( .A1(ymem_data1[42]), .A2(n3289), .B1(n3202), .B2(
        U72_DATA1_42), .C1(ymem_data1[106]), .C2(n3288), .ZN(n1880) );
  AOI21_X2 U1778 ( .B1(n1882), .B2(n1883), .A(n3286), .ZN(n1881) );
  AOI21_X2 U1780 ( .B1(n1872), .B2(n1873), .A(n3300), .ZN(U94_Z_43) );
  AOI222_X1 U1782 ( .A1(ymem_data1[43]), .A2(n3289), .B1(n3202), .B2(
        U72_DATA1_43), .C1(ymem_data1[107]), .C2(n3288), .ZN(n1873) );
  AOI21_X2 U1784 ( .B1(n1875), .B2(n1876), .A(n3286), .ZN(n1874) );
  AOI21_X2 U1787 ( .B1(n1865), .B2(n1866), .A(n3300), .ZN(U94_Z_44) );
  AOI222_X1 U1789 ( .A1(ymem_data1[44]), .A2(n628), .B1(n3202), .B2(
        U72_DATA1_44), .C1(ymem_data1[108]), .C2(n3288), .ZN(n1866) );
  AOI21_X2 U1791 ( .B1(n1868), .B2(n1869), .A(n3286), .ZN(n1867) );
  AOI21_X2 U1793 ( .B1(n1858), .B2(n1859), .A(n3300), .ZN(U94_Z_45) );
  AOI222_X1 U1794 ( .A1(ymem_data1[45]), .A2(n628), .B1(n3202), .B2(
        U72_DATA1_45), .C1(ymem_data1[109]), .C2(n3288), .ZN(n1859) );
  AOI21_X2 U1795 ( .B1(n1861), .B2(n1862), .A(n3286), .ZN(n1860) );
  AOI21_X2 U1907 ( .B1(n1851), .B2(n1852), .A(n3300), .ZN(U94_Z_46) );
  AOI222_X1 U1909 ( .A1(ymem_data1[46]), .A2(n3289), .B1(n3202), .B2(
        U72_DATA1_46), .C1(ymem_data1[110]), .C2(n3288), .ZN(n1852) );
  AOI21_X2 U1911 ( .B1(n1854), .B2(n1855), .A(n3286), .ZN(n1853) );
  AOI21_X2 U1916 ( .B1(n1844), .B2(n1845), .A(n3300), .ZN(U94_Z_47) );
  AOI222_X1 U1919 ( .A1(ymem_data1[47]), .A2(n628), .B1(n3202), .B2(
        U72_DATA1_47), .C1(ymem_data1[111]), .C2(n3288), .ZN(n1845) );
  AOI21_X2 U1922 ( .B1(n1847), .B2(n1848), .A(n3286), .ZN(n1846) );
  AOI22_X2 U1925 ( .A1(ymem_data2[52]), .A2(n2472), .B1(ymem_data1[180]), .B2(
        n3287), .ZN(n2484) );
  AOI22_X2 U1929 ( .A1(ymem_data2[56]), .A2(n2472), .B1(ymem_data1[184]), .B2(
        n3287), .ZN(n2492) );
  AOI22_X2 U1932 ( .A1(ymem_data2[60]), .A2(n2472), .B1(ymem_data1[188]), .B2(
        n3287), .ZN(n2500) );
  AOI22_X2 U1935 ( .A1(ymem_data2[59]), .A2(n2472), .B1(ymem_data1[187]), .B2(
        n3287), .ZN(n2489) );
  NAND3_X2 U1938 ( .A1(n152), .A2(n149), .A3(n[2371]), .ZN(n2156) );
  AOI22_X2 U1942 ( .A1(ymem_data2[53]), .A2(n2472), .B1(ymem_data1[181]), .B2(
        n3287), .ZN(n2483) );
  AOI22_X2 U1945 ( .A1(ymem_data2[57]), .A2(n2472), .B1(ymem_data1[185]), .B2(
        n3287), .ZN(n2491) );
  AOI22_X2 U1948 ( .A1(ymem_data2[61]), .A2(n2472), .B1(ymem_data1[189]), .B2(
        n3287), .ZN(n2499) );
  AOI22_X2 U1951 ( .A1(ymem_data2[58]), .A2(n2472), .B1(ymem_data1[186]), .B2(
        n3287), .ZN(n2490) );
  AOI22_X2 U1955 ( .A1(ymem_data2[62]), .A2(n2472), .B1(ymem_data1[190]), .B2(
        n3287), .ZN(n2498) );
  AOI22_X2 U1958 ( .A1(ymem_data1[248]), .A2(n128), .B1(ymem_data1[249]), .B2(
        n127), .ZN(n2563) );
  INV_X4 U1964 ( .A(n715), .ZN(n3287) );
  INV_X4 U1965 ( .A(n1811), .ZN(n3226) );
  OAI222_X2 U1970 ( .A1(n2246), .A2(n384), .B1(n2247), .B2(n256), .C1(n715), 
        .C2(n576), .ZN(n2250) );
  OAI222_X2 U1976 ( .A1(n2246), .A2(n385), .B1(n2247), .B2(n257), .C1(n715), 
        .C2(n577), .ZN(n2252) );
  OAI222_X2 U1986 ( .A1(n2246), .A2(n386), .B1(n2247), .B2(n258), .C1(n715), 
        .C2(n578), .ZN(n2254) );
  AOI21_X2 U1989 ( .B1(chng_row[15]), .B2(n113), .A(n2227), .ZN(n2283) );
  OAI222_X2 U1991 ( .A1(n2246), .A2(n371), .B1(n2247), .B2(n243), .C1(n715), 
        .C2(n563), .ZN(n2284) );
  AOI21_X2 U1993 ( .B1(chng_row[14]), .B2(n113), .A(n2229), .ZN(n2285) );
  OAI222_X2 U1996 ( .A1(n2246), .A2(n372), .B1(n2247), .B2(n244), .C1(n715), 
        .C2(n564), .ZN(n2286) );
  AOI22_X2 U2000 ( .A1(ymem_data1[0]), .A2(n3295), .B1(ymem_data2[192]), .B2(
        n3298), .ZN(n871) );
  AOI22_X2 U2003 ( .A1(ymem_data1[34]), .A2(n3295), .B1(ymem_data2[226]), .B2(
        n3298), .ZN(n1517) );
  AOI22_X2 U2006 ( .A1(ymem_data1[32]), .A2(n3295), .B1(ymem_data2[224]), .B2(
        n3298), .ZN(n1479) );
  AOI22_X2 U2009 ( .A1(ymem_data1[31]), .A2(n3295), .B1(ymem_data2[223]), .B2(
        n3298), .ZN(n1460) );
  AOI22_X2 U2013 ( .A1(ymem_data1[30]), .A2(n3295), .B1(ymem_data2[222]), .B2(
        n3298), .ZN(n1441) );
  AOI22_X2 U2016 ( .A1(ymem_data1[29]), .A2(n3295), .B1(ymem_data2[221]), .B2(
        n3298), .ZN(n1422) );
  AOI22_X2 U2019 ( .A1(ymem_data1[28]), .A2(n3295), .B1(ymem_data2[220]), .B2(
        n3298), .ZN(n1403) );
  AOI22_X2 U2021 ( .A1(ymem_data1[27]), .A2(n3295), .B1(ymem_data2[219]), .B2(
        n3298), .ZN(n1384) );
  AOI22_X2 U2069 ( .A1(ymem_data1[26]), .A2(n3295), .B1(ymem_data2[218]), .B2(
        n3298), .ZN(n1365) );
  AOI22_X2 U2072 ( .A1(ymem_data1[25]), .A2(n3295), .B1(ymem_data2[217]), .B2(
        n3298), .ZN(n1346) );
  AOI22_X2 U2075 ( .A1(ymem_data1[24]), .A2(n3295), .B1(ymem_data2[216]), .B2(
        n3298), .ZN(n1327) );
  AOI22_X2 U2078 ( .A1(ymem_data1[23]), .A2(n3295), .B1(ymem_data2[215]), .B2(
        n3298), .ZN(n1308) );
  AOI22_X2 U2082 ( .A1(ymem_data1[22]), .A2(n3295), .B1(ymem_data2[214]), .B2(
        n3298), .ZN(n1289) );
  AOI22_X2 U2092 ( .A1(ymem_data1[21]), .A2(n3295), .B1(ymem_data2[213]), .B2(
        n3298), .ZN(n1270) );
  AOI22_X2 U2094 ( .A1(ymem_data1[20]), .A2(n3295), .B1(ymem_data2[212]), .B2(
        n3298), .ZN(n1251) );
  AOI22_X2 U2097 ( .A1(ymem_data1[19]), .A2(n3295), .B1(ymem_data2[211]), .B2(
        n3298), .ZN(n1232) );
  AOI22_X2 U2099 ( .A1(ymem_data1[17]), .A2(n3295), .B1(ymem_data2[209]), .B2(
        n3298), .ZN(n1194) );
  AOI22_X2 U2108 ( .A1(ymem_data1[16]), .A2(n3295), .B1(ymem_data2[208]), .B2(
        n3298), .ZN(n1175) );
  AOI22_X2 U2125 ( .A1(ymem_data1[15]), .A2(n3295), .B1(ymem_data2[207]), .B2(
        n3298), .ZN(n1156) );
  AOI22_X2 U2127 ( .A1(ymem_data1[14]), .A2(n3295), .B1(ymem_data2[206]), .B2(
        n3298), .ZN(n1137) );
  AOI22_X2 U2145 ( .A1(ymem_data1[13]), .A2(n3295), .B1(ymem_data2[205]), .B2(
        n3298), .ZN(n1118) );
  AOI22_X2 U2156 ( .A1(ymem_data1[12]), .A2(n3295), .B1(ymem_data2[204]), .B2(
        n3298), .ZN(n1099) );
  AOI22_X2 U2157 ( .A1(ymem_data1[11]), .A2(n3295), .B1(ymem_data2[203]), .B2(
        n3298), .ZN(n1080) );
  AOI22_X2 U2159 ( .A1(ymem_data1[35]), .A2(n3295), .B1(ymem_data2[227]), .B2(
        n3298), .ZN(n1536) );
  AOI22_X2 U2161 ( .A1(ymem_data1[33]), .A2(n3295), .B1(ymem_data2[225]), .B2(
        n3298), .ZN(n1498) );
  AOI22_X2 U2166 ( .A1(ymem_data1[18]), .A2(n3295), .B1(ymem_data2[210]), .B2(
        n3298), .ZN(n1213) );
  AOI22_X2 U2167 ( .A1(ymem_data1[10]), .A2(n3295), .B1(ymem_data2[202]), .B2(
        n3298), .ZN(n1061) );
  AOI22_X2 U2172 ( .A1(ymem_data1[9]), .A2(n3295), .B1(ymem_data2[201]), .B2(
        n3298), .ZN(n1042) );
  AOI22_X2 U2176 ( .A1(ymem_data1[8]), .A2(n3295), .B1(ymem_data2[200]), .B2(
        n3298), .ZN(n1023) );
  AOI22_X2 U2183 ( .A1(ymem_data1[7]), .A2(n3295), .B1(ymem_data2[199]), .B2(
        n3298), .ZN(n1004) );
  AOI22_X2 U2185 ( .A1(ymem_data1[6]), .A2(n3295), .B1(ymem_data2[198]), .B2(
        n3298), .ZN(n985) );
  AOI22_X2 U2193 ( .A1(ymem_data1[5]), .A2(n3295), .B1(ymem_data2[197]), .B2(
        n3298), .ZN(n966) );
  AOI22_X2 U2195 ( .A1(ymem_data1[4]), .A2(n3295), .B1(ymem_data2[196]), .B2(
        n3298), .ZN(n947) );
  AOI22_X2 U2196 ( .A1(ymem_data1[3]), .A2(n3295), .B1(ymem_data2[195]), .B2(
        n3298), .ZN(n928) );
  AOI22_X2 U2197 ( .A1(ymem_data1[2]), .A2(n3295), .B1(ymem_data2[194]), .B2(
        n3298), .ZN(n909) );
  AOI22_X2 U2199 ( .A1(ymem_data1[1]), .A2(n3295), .B1(ymem_data2[193]), .B2(
        n3298), .ZN(n890) );
  OAI21_X2 U2200 ( .B1(n3301), .B2(n1790), .A(n1791), .ZN(U95_Z_1) );
  AOI22_X2 U2201 ( .A1(n150), .A2(chng_col[6]), .B1(n3291), .B2(chng_row[6]), 
        .ZN(n2542) );
  AOI22_X2 U2202 ( .A1(n150), .A2(chng_col[5]), .B1(n3291), .B2(chng_row[5]), 
        .ZN(n2539) );
  AOI22_X2 U2203 ( .A1(n150), .A2(chng_col[7]), .B1(n3291), .B2(chng_row[7]), 
        .ZN(n2545) );
  AOI22_X2 U2678 ( .A1(n150), .A2(chng_col[0]), .B1(n3291), .B2(chng_row[0]), 
        .ZN(n2525) );
  AOI22_X2 U2680 ( .A1(n150), .A2(chng_col[1]), .B1(n3291), .B2(chng_row[1]), 
        .ZN(n2528) );
  AOI22_X2 U2684 ( .A1(n150), .A2(chng_col[4]), .B1(n3291), .B2(chng_row[4]), 
        .ZN(n2536) );
  AOI22_X2 U2733 ( .A1(chng_row[2]), .A2(n2301), .B1(chng_col[2]), .B2(n2302), 
        .ZN(n2303) );
  AOI22_X2 U2735 ( .A1(chng_row[1]), .A2(n2301), .B1(chng_col[1]), .B2(n2302), 
        .ZN(n2304) );
  AOI22_X2 U2736 ( .A1(chng_row[0]), .A2(n2301), .B1(chng_col[0]), .B2(n2302), 
        .ZN(n2305) );
  AOI22_X2 U2738 ( .A1(chng_row[3]), .A2(n2301), .B1(chng_col[3]), .B2(n2302), 
        .ZN(n2300) );
  AOI22_X2 U2742 ( .A1(chng_row[7]), .A2(n2301), .B1(chng_col[7]), .B2(n2302), 
        .ZN(n2310) );
  AOI22_X2 U2743 ( .A1(chng_row[5]), .A2(n2301), .B1(chng_col[5]), .B2(n2302), 
        .ZN(n2312) );
  AOI22_X2 U2744 ( .A1(chng_row[4]), .A2(n2301), .B1(chng_col[4]), .B2(n2302), 
        .ZN(n2313) );
  AOI22_X2 U2745 ( .A1(chng_row[11]), .A2(n2301), .B1(chng_col[11]), .B2(n2302), .ZN(n2318) );
  AOI22_X2 U2746 ( .A1(chng_row[9]), .A2(n2301), .B1(chng_col[9]), .B2(n2302), 
        .ZN(n2320) );
  AOI22_X2 U2747 ( .A1(chng_row[8]), .A2(n2301), .B1(chng_col[8]), .B2(n2302), 
        .ZN(n2321) );
  AOI22_X2 U2748 ( .A1(chng_row[15]), .A2(n2301), .B1(chng_col[15]), .B2(n2302), .ZN(n2326) );
  AOI22_X2 U2749 ( .A1(chng_row[13]), .A2(n2301), .B1(chng_col[13]), .B2(n2302), .ZN(n2328) );
  AOI22_X2 U2750 ( .A1(chng_row[12]), .A2(n2301), .B1(chng_col[12]), .B2(n2302), .ZN(n2329) );
  AOI22_X2 U2751 ( .A1(ymem_data1[114]), .A2(n3291), .B1(ymem_data1[50]), .B2(
        n150), .ZN(n2612) );
  AOI22_X2 U2752 ( .A1(ymem_data1[46]), .A2(n3295), .B1(ymem_data2[238]), .B2(
        n3298), .ZN(n1745) );
  AOI22_X2 U2753 ( .A1(ymem_data1[45]), .A2(n3295), .B1(ymem_data2[237]), .B2(
        n3298), .ZN(n1726) );
  AOI22_X2 U2754 ( .A1(ymem_data1[44]), .A2(n3295), .B1(ymem_data2[236]), .B2(
        n3298), .ZN(n1707) );
  AOI22_X2 U2755 ( .A1(ymem_data1[43]), .A2(n3295), .B1(ymem_data2[235]), .B2(
        n3298), .ZN(n1688) );
  AOI22_X2 U2756 ( .A1(ymem_data1[42]), .A2(n3295), .B1(ymem_data2[234]), .B2(
        n3298), .ZN(n1669) );
  AOI22_X2 U2757 ( .A1(ymem_data1[41]), .A2(n3295), .B1(ymem_data2[233]), .B2(
        n3298), .ZN(n1650) );
  AOI22_X2 U2758 ( .A1(ymem_data1[40]), .A2(n3295), .B1(ymem_data2[232]), .B2(
        n3298), .ZN(n1631) );
  AOI22_X2 U2759 ( .A1(ymem_data1[39]), .A2(n3295), .B1(ymem_data2[231]), .B2(
        n3298), .ZN(n1612) );
  AOI22_X2 U2760 ( .A1(ymem_data1[38]), .A2(n3295), .B1(ymem_data2[230]), .B2(
        n3298), .ZN(n1593) );
  AOI22_X2 U2761 ( .A1(ymem_data1[37]), .A2(n3295), .B1(ymem_data2[229]), .B2(
        n3298), .ZN(n1574) );
  AOI22_X2 U2762 ( .A1(ymem_data1[36]), .A2(n3295), .B1(ymem_data2[228]), .B2(
        n3298), .ZN(n1555) );
  AOI22_X2 U2763 ( .A1(ymem_data1[47]), .A2(n3295), .B1(ymem_data2[239]), .B2(
        n3298), .ZN(n1779) );
  AOI22_X2 U2764 ( .A1(n8), .A2(n767), .B1(op_oneHotNonDiag[0]), .B2(n7), .ZN(
        n766) );
  AOI222_X1 U2765 ( .A1(n736), .A2(n3279), .B1(n117), .B2(n91), .C1(n139), 
        .C2(n90), .ZN(n769) );
  AOI22_X2 U2766 ( .A1(chng_row[6]), .A2(n2301), .B1(chng_col[6]), .B2(n2302), 
        .ZN(n2311) );
  AOI22_X2 U2767 ( .A1(chng_row[10]), .A2(n2301), .B1(chng_col[10]), .B2(n2302), .ZN(n2319) );
  AOI22_X2 U2768 ( .A1(chng_row[14]), .A2(n2301), .B1(chng_col[14]), .B2(n2302), .ZN(n2327) );
  AOI21_X2 U2769 ( .B1(chng_row[2]), .B2(n113), .A(n2193), .ZN(n2249) );
  AOI21_X2 U2770 ( .B1(chng_row[1]), .B2(n113), .A(n2195), .ZN(n2251) );
  AOI21_X2 U2771 ( .B1(chng_row[0]), .B2(n113), .A(n2197), .ZN(n2253) );
  AOI21_X2 U2772 ( .B1(chng_row[4]), .B2(n113), .A(n2209), .ZN(n2265) );
  OAI222_X2 U2773 ( .A1(n2246), .A2(n382), .B1(n2247), .B2(n254), .C1(n715), 
        .C2(n574), .ZN(n2266) );
  AOI21_X2 U2774 ( .B1(chng_row[8]), .B2(n113), .A(n2221), .ZN(n2277) );
  OAI222_X2 U2775 ( .A1(n2246), .A2(n378), .B1(n2247), .B2(n250), .C1(n715), 
        .C2(n570), .ZN(n2278) );
  AOI21_X2 U2776 ( .B1(chng_row[12]), .B2(n113), .A(n2233), .ZN(n2289) );
  OAI222_X2 U2777 ( .A1(n2246), .A2(n374), .B1(n2247), .B2(n246), .C1(n715), 
        .C2(n566), .ZN(n2290) );
  AOI21_X2 U2778 ( .B1(chng_row[3]), .B2(n113), .A(n2190), .ZN(n2244) );
  OAI222_X2 U2779 ( .A1(n2246), .A2(n383), .B1(n2247), .B2(n255), .C1(n3286), 
        .C2(n575), .ZN(n2245) );
  AOI21_X2 U2780 ( .B1(chng_row[7]), .B2(n113), .A(n2203), .ZN(n2259) );
  OAI222_X2 U2781 ( .A1(n2246), .A2(n379), .B1(n2247), .B2(n251), .C1(n3286), 
        .C2(n571), .ZN(n2260) );
  AOI21_X2 U2782 ( .B1(chng_row[11]), .B2(n113), .A(n2215), .ZN(n2271) );
  OAI222_X2 U2783 ( .A1(n2246), .A2(n375), .B1(n2247), .B2(n247), .C1(n715), 
        .C2(n567), .ZN(n2272) );
  AOI21_X2 U2784 ( .B1(chng_row[5]), .B2(n113), .A(n2207), .ZN(n2263) );
  OAI222_X2 U2785 ( .A1(n2246), .A2(n381), .B1(n2247), .B2(n253), .C1(n715), 
        .C2(n573), .ZN(n2264) );
  AOI21_X2 U2786 ( .B1(chng_row[9]), .B2(n113), .A(n2219), .ZN(n2275) );
  OAI222_X2 U2787 ( .A1(n2246), .A2(n377), .B1(n2247), .B2(n249), .C1(n715), 
        .C2(n569), .ZN(n2276) );
  AOI21_X2 U2788 ( .B1(chng_row[13]), .B2(n113), .A(n2231), .ZN(n2287) );
  OAI222_X2 U2789 ( .A1(n2246), .A2(n373), .B1(n2247), .B2(n245), .C1(n715), 
        .C2(n565), .ZN(n2288) );
  AOI21_X2 U2790 ( .B1(chng_row[6]), .B2(n113), .A(n2205), .ZN(n2261) );
  OAI222_X2 U2791 ( .A1(n2246), .A2(n380), .B1(n2247), .B2(n252), .C1(n715), 
        .C2(n572), .ZN(n2262) );
  AOI21_X2 U2792 ( .B1(chng_row[10]), .B2(n113), .A(n2217), .ZN(n2273) );
  OAI222_X2 U2793 ( .A1(n2246), .A2(n376), .B1(n2247), .B2(n248), .C1(n715), 
        .C2(n568), .ZN(n2274) );
  OAI21_X2 U2794 ( .B1(n806), .B2(n786), .A(n807), .ZN(n2629) );
  OAI21_X2 U2795 ( .B1(n3301), .B2(n1793), .A(n134), .ZN(U95_Z_0) );
  INV_X4 U2797 ( .A(n1815), .ZN(n3222) );
  AOI22_X2 U2798 ( .A1(ymem_data1[115]), .A2(n3291), .B1(ymem_data1[51]), .B2(
        n150), .ZN(n2613) );
  OAI21_X2 U2799 ( .B1(n820), .B2(n821), .A(n8), .ZN(n819) );
  OAI21_X2 U2800 ( .B1(n3214), .B2(n629), .A(n630), .ZN(n2614) );
  AOI22_X2 U2801 ( .A1(n73), .A2(n628), .B1(op_oneHotDiag[0]), .B2(n72), .ZN(
        n627) );
  AOI21_X2 U2802 ( .B1(n[2370]), .B2(n133), .A(n828), .ZN(n1772) );
  OAI21_X2 U2803 ( .B1(n2151), .B2(n765), .A(reset), .ZN(n2150) );
  INV_X4 U2804 ( .A(n3215), .ZN(n3221) );
  AND2_X4 U2805 ( .A1(n2387), .A2(n3278), .ZN(n2473) );
  AND2_X4 U2806 ( .A1(n3205), .A2(n2387), .ZN(n2340) );
  NAND3_X2 U2807 ( .A1(n[2370]), .A2(n151), .A3(n[2372]), .ZN(n3218) );
  NAND3_X2 U2808 ( .A1(n[2370]), .A2(n151), .A3(n[2372]), .ZN(n3219) );
  AND3_X4 U2809 ( .A1(n717), .A2(n795), .A3(n2235), .ZN(n2192) );
  NAND3_X1 U3 ( .A1(n829), .A2(n3221), .A3(n831), .ZN(n764) );
  INV_X2 U9 ( .A(n854), .ZN(n3260) );
  INV_X1 U14 ( .A(n3197), .ZN(n3302) );
  INV_X8 U84 ( .A(n3302), .ZN(n3303) );
  NAND2_X2 U103 ( .A1(n752), .A2(n3259), .ZN(n3197) );
  INV_X8 U109 ( .A(n3267), .ZN(n3266) );
  INV_X8 U144 ( .A(n1780), .ZN(n3298) );
  AOI221_X1 U156 ( .B1(ymem_data1[219]), .B2(n3283), .C1(ymem_data1[155]), 
        .C2(n782), .A(n2000), .ZN(n1998) );
  AOI221_X1 U163 ( .B1(ymem_data1[194]), .B2(n3283), .C1(ymem_data1[130]), 
        .C2(n782), .A(n2056), .ZN(n2054) );
  AOI221_X1 U172 ( .B1(ymem_data1[207]), .B2(n3283), .C1(ymem_data1[143]), 
        .C2(n782), .A(n2091), .ZN(n2089) );
  AOI221_X1 U239 ( .B1(ymem_data1[206]), .B2(n3283), .C1(ymem_data1[142]), 
        .C2(n782), .A(n2098), .ZN(n2096) );
  AOI221_X1 U246 ( .B1(ymem_data2[135]), .B2(n3270), .C1(ymem_data2[199]), 
        .C2(n849), .A(n997), .ZN(n996) );
  AOI221_X1 U276 ( .B1(ymem_data2[138]), .B2(n3271), .C1(ymem_data2[202]), 
        .C2(n849), .A(n1054), .ZN(n1053) );
  AOI221_X1 U293 ( .B1(ymem_data2[140]), .B2(n3271), .C1(ymem_data2[204]), 
        .C2(n849), .A(n1092), .ZN(n1091) );
  AOI221_X1 U316 ( .B1(ymem_data2[141]), .B2(n3271), .C1(ymem_data2[205]), 
        .C2(n849), .A(n1111), .ZN(n1110) );
  AOI221_X1 U353 ( .B1(n3234), .B2(ymem_data2[204]), .C1(n1807), .C2(
        ymem_data1[12]), .A(n2115), .ZN(n2114) );
  AOI221_X1 U391 ( .B1(n3235), .B2(ymem_data2[203]), .C1(n1807), .C2(
        ymem_data1[11]), .A(n2122), .ZN(n2121) );
  AOI221_X1 U393 ( .B1(n3234), .B2(ymem_data2[202]), .C1(n1807), .C2(
        ymem_data1[10]), .A(n2129), .ZN(n2128) );
  AOI221_X1 U413 ( .B1(n3235), .B2(ymem_data2[193]), .C1(n1807), .C2(
        ymem_data1[1]), .A(n2136), .ZN(n2135) );
  AOI21_X1 U419 ( .B1(n2001), .B2(n2002), .A(n715), .ZN(n2000) );
  AOI21_X1 U423 ( .B1(n1987), .B2(n1988), .A(n715), .ZN(n1986) );
  AOI21_X1 U439 ( .B1(n1966), .B2(n1967), .A(n715), .ZN(n1965) );
  AOI21_X1 U443 ( .B1(n2029), .B2(n2030), .A(n715), .ZN(n2028) );
  AOI21_X1 U459 ( .B1(n2015), .B2(n2016), .A(n715), .ZN(n2014) );
  OAI222_X1 U584 ( .A1(n829), .A2(n1799), .B1(n2), .B2(n715), .C1(
        yMemDataReadyNextCycle), .C2(n3221), .ZN(n1795) );
  OAI22_X1 U586 ( .A1(n794), .A2(n442), .B1(n2192), .B2(n314), .ZN(n2222) );
  OAI22_X1 U596 ( .A1(n794), .A2(n446), .B1(n2192), .B2(n318), .ZN(n2210) );
  OAI22_X1 U606 ( .A1(n794), .A2(n437), .B1(n2192), .B2(n309), .ZN(n2232) );
  OAI22_X1 U612 ( .A1(n450), .A2(n794), .B1(n2192), .B2(n322), .ZN(n2198) );
  OAI222_X1 U616 ( .A1(n554), .A2(n3230), .B1(n618), .B2(n1810), .C1(n490), 
        .C2(n1811), .ZN(n1821) );
  OAI222_X1 U636 ( .A1(n553), .A2(n3231), .B1(n617), .B2(n1810), .C1(n489), 
        .C2(n1811), .ZN(n1808) );
  OAI222_X1 U639 ( .A1(n532), .A2(n3230), .B1(n596), .B2(n1810), .C1(n468), 
        .C2(n3227), .ZN(n1975) );
  OAI222_X1 U646 ( .A1(n546), .A2(n3230), .B1(n610), .B2(n1810), .C1(n482), 
        .C2(n1811), .ZN(n2087) );
  OAI222_X1 U656 ( .A1(n544), .A2(n3230), .B1(n608), .B2(n1810), .C1(n480), 
        .C2(n1811), .ZN(n2073) );
  OAI221_X1 U659 ( .B1(n3248), .B2(n262), .C1(n870), .C2(n326), .A(n1707), 
        .ZN(n1705) );
  OAI221_X1 U679 ( .B1(n3248), .B2(n260), .C1(n870), .C2(n324), .A(n1745), 
        .ZN(n1743) );
  OAI221_X1 U739 ( .B1(n306), .B2(n3248), .C1(n870), .C2(n370), .A(n871), .ZN(
        n867) );
  OAI221_X1 U759 ( .B1(n3249), .B2(n293), .C1(n870), .C2(n357), .A(n1118), 
        .ZN(n1116) );
  OAI221_X1 U779 ( .B1(n3249), .B2(n292), .C1(n870), .C2(n356), .A(n1137), 
        .ZN(n1135) );
  OAI22_X1 U839 ( .A1(n777), .A2(n778), .B1(n779), .B2(n3286), .ZN(n772) );
  OAI22_X1 U991 ( .A1(n3307), .A2(n326), .B1(n778), .B2(n390), .ZN(n1697) );
  OAI22_X1 U1011 ( .A1(n3307), .A2(n327), .B1(n778), .B2(n391), .ZN(n1678) );
  OAI22_X1 U1031 ( .A1(n3307), .A2(n328), .B1(n778), .B2(n392), .ZN(n1659) );
  OAI22_X1 U1043 ( .A1(n3307), .A2(n358), .B1(n778), .B2(n422), .ZN(n1089) );
  INV_X1 U1083 ( .A(n3196), .ZN(n3304) );
  INV_X8 U1390 ( .A(n3304), .ZN(n3305) );
  NAND2_X2 U1454 ( .A1(n751), .A2(n3259), .ZN(n3196) );
  OAI22_X1 U1494 ( .A1(n294), .A2(n3198), .B1(n358), .B2(n1815), .ZN(n2116) );
  OAI22_X1 U1499 ( .A1(n295), .A2(n3198), .B1(n359), .B2(n1815), .ZN(n2123) );
  OAI22_X1 U1502 ( .A1(n296), .A2(n3198), .B1(n360), .B2(n1815), .ZN(n2130) );
  OAI22_X1 U1520 ( .A1(n305), .A2(n3198), .B1(n369), .B2(n1815), .ZN(n2137) );
  OAI22_X1 U1523 ( .A1(n306), .A2(n3198), .B1(n370), .B2(n1815), .ZN(n2148) );
  OAI22_X1 U1528 ( .A1(n291), .A2(n3198), .B1(n355), .B2(n1815), .ZN(n2095) );
  OAI22_X1 U1531 ( .A1(n862), .A2(n339), .B1(n3248), .B2(n275), .ZN(n1457) );
  OAI22_X1 U1536 ( .A1(n862), .A2(n341), .B1(n3249), .B2(n277), .ZN(n1419) );
  OAI22_X1 U1539 ( .A1(n862), .A2(n340), .B1(n3249), .B2(n276), .ZN(n1438) );
  OAI22_X1 U1544 ( .A1(n862), .A2(n357), .B1(n3249), .B2(n293), .ZN(n1115) );
  OAI22_X1 U1547 ( .A1(n862), .A2(n356), .B1(n3249), .B2(n292), .ZN(n1134) );
  OAI22_X1 U1558 ( .A1(n862), .A2(n355), .B1(n3249), .B2(n291), .ZN(n1153) );
  OAI22_X1 U1577 ( .A1(n862), .A2(n336), .B1(n3249), .B2(n272), .ZN(n1514) );
  OAI22_X1 U1586 ( .A1(n862), .A2(n366), .B1(n863), .B2(n302), .ZN(n944) );
  OAI22_X1 U1638 ( .A1(n862), .A2(n346), .B1(n863), .B2(n282), .ZN(n1324) );
  OAI22_X1 U1654 ( .A1(n862), .A2(n345), .B1(n863), .B2(n281), .ZN(n1343) );
  OAI22_X1 U1663 ( .A1(n862), .A2(n344), .B1(n863), .B2(n280), .ZN(n1362) );
  OAI22_X1 U1672 ( .A1(n856), .A2(n236), .B1(n3255), .B2(n300), .ZN(n979) );
  OAI22_X1 U1679 ( .A1(n856), .A2(n234), .B1(n3255), .B2(n298), .ZN(n1017) );
  OAI22_X1 U1692 ( .A1(n856), .A2(n220), .B1(n3255), .B2(n284), .ZN(n1283) );
  OAI22_X1 U1705 ( .A1(n856), .A2(n219), .B1(n3255), .B2(n283), .ZN(n1302) );
  OAI22_X1 U1961 ( .A1(n856), .A2(n218), .B1(n3255), .B2(n282), .ZN(n1321) );
  OAI22_X1 U2796 ( .A1(n856), .A2(n217), .B1(n3255), .B2(n281), .ZN(n1340) );
  OAI22_X1 U2810 ( .A1(n856), .A2(n242), .B1(n3255), .B2(n306), .ZN(n855) );
  INV_X1 U2811 ( .A(n3199), .ZN(n3306) );
  INV_X8 U2812 ( .A(n3306), .ZN(n3307) );
  NAND2_X2 U2813 ( .A1(n112), .A2(n3259), .ZN(n3199) );
  INV_X8 U2814 ( .A(n1768), .ZN(n3299) );
  INV_X1 U2815 ( .A(n834), .ZN(n3308) );
  INV_X8 U2816 ( .A(n3308), .ZN(n3309) );
  INV_X8 U2817 ( .A(n3287), .ZN(n3286) );
endmodule


module getYMatAddress ( readEnable, gYMA_row, gYMA_readData, gYMA_row_addr1 );
  input [15:0] gYMA_row;
  input [255:0] gYMA_readData;
  output [10:0] gYMA_row_addr1;
  input readEnable;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;

  AND4_X2 U3 ( .A1(n6), .A2(n7), .A3(n8), .A4(n9), .ZN(n5) );
  AND4_X2 U8 ( .A1(n18), .A2(n19), .A3(n20), .A4(n21), .ZN(n4) );
  AND4_X2 U14 ( .A1(n32), .A2(n33), .A3(n34), .A4(n35), .ZN(n31) );
  AND4_X2 U19 ( .A1(n36), .A2(n37), .A3(n38), .A4(n39), .ZN(n30) );
  AND4_X2 U25 ( .A1(n42), .A2(n43), .A3(n44), .A4(n45), .ZN(n41) );
  AND4_X2 U30 ( .A1(n46), .A2(n47), .A3(n48), .A4(n49), .ZN(n40) );
  AND4_X2 U36 ( .A1(n52), .A2(n53), .A3(n54), .A4(n55), .ZN(n51) );
  AND4_X2 U41 ( .A1(n56), .A2(n57), .A3(n58), .A4(n59), .ZN(n50) );
  AND4_X2 U47 ( .A1(n62), .A2(n63), .A3(n64), .A4(n65), .ZN(n61) );
  AND4_X2 U52 ( .A1(n66), .A2(n67), .A3(n68), .A4(n69), .ZN(n60) );
  AND4_X2 U58 ( .A1(n72), .A2(n73), .A3(n74), .A4(n75), .ZN(n71) );
  AND4_X2 U63 ( .A1(n76), .A2(n77), .A3(n78), .A4(n79), .ZN(n70) );
  AND4_X2 U69 ( .A1(n82), .A2(n83), .A3(n84), .A4(n85), .ZN(n81) );
  AND4_X2 U74 ( .A1(n86), .A2(n87), .A3(n88), .A4(n89), .ZN(n80) );
  AND4_X2 U80 ( .A1(n92), .A2(n93), .A3(n94), .A4(n95), .ZN(n91) );
  AND4_X2 U85 ( .A1(n96), .A2(n97), .A3(n98), .A4(n99), .ZN(n90) );
  AND4_X2 U91 ( .A1(n102), .A2(n103), .A3(n104), .A4(n105), .ZN(n101) );
  AND4_X2 U96 ( .A1(n106), .A2(n107), .A3(n108), .A4(n109), .ZN(n100) );
  AND4_X2 U102 ( .A1(n112), .A2(n113), .A3(n114), .A4(n115), .ZN(n111) );
  AND4_X2 U107 ( .A1(n122), .A2(n123), .A3(n124), .A4(n125), .ZN(n110) );
  NOR2_X2 U111 ( .A1(n2), .A2(gYMA_row[2]), .ZN(n120) );
  NOR2_X2 U113 ( .A1(gYMA_row[3]), .A2(gYMA_row[0]), .ZN(n126) );
  NOR2_X2 U114 ( .A1(gYMA_row[2]), .A2(gYMA_row[1]), .ZN(n121) );
  NOR2_X2 U115 ( .A1(n3), .A2(gYMA_row[3]), .ZN(n127) );
  INV_X4 U117 ( .A(gYMA_row[1]), .ZN(n2) );
  INV_X4 U118 ( .A(gYMA_row[0]), .ZN(n3) );
  AND2_X1 U126 ( .A1(gYMA_row[3]), .A2(n3), .ZN(n116) );
  AND2_X1 U128 ( .A1(gYMA_row[3]), .A2(gYMA_row[0]), .ZN(n118) );
  AND2_X1 U131 ( .A1(gYMA_row[2]), .A2(gYMA_row[1]), .ZN(n117) );
  AND2_X1 U134 ( .A1(gYMA_row[2]), .A2(n2), .ZN(n119) );
  INV_X4 U2 ( .A(1'b1), .ZN(gYMA_row_addr1[10]) );
  AOI21_X2 U5 ( .B1(n100), .B2(n101), .A(n1), .ZN(gYMA_row_addr1[1]) );
  AOI22_X2 U6 ( .A1(gYMA_readData[225]), .A2(n28), .B1(gYMA_readData[241]), 
        .B2(n29), .ZN(n106) );
  AOI21_X2 U7 ( .B1(n110), .B2(n111), .A(n1), .ZN(gYMA_row_addr1[0]) );
  AOI22_X2 U9 ( .A1(gYMA_readData[224]), .A2(n28), .B1(gYMA_readData[240]), 
        .B2(n29), .ZN(n122) );
  AOI21_X2 U10 ( .B1(n80), .B2(n81), .A(n1), .ZN(gYMA_row_addr1[3]) );
  AOI22_X2 U11 ( .A1(gYMA_readData[227]), .A2(n28), .B1(gYMA_readData[243]), 
        .B2(n29), .ZN(n86) );
  AOI21_X2 U12 ( .B1(n90), .B2(n91), .A(n1), .ZN(gYMA_row_addr1[2]) );
  AOI22_X2 U13 ( .A1(gYMA_readData[226]), .A2(n28), .B1(gYMA_readData[242]), 
        .B2(n29), .ZN(n96) );
  AOI22_X2 U15 ( .A1(gYMA_readData[64]), .A2(n14), .B1(gYMA_readData[80]), 
        .B2(n15), .ZN(n113) );
  AOI22_X2 U16 ( .A1(gYMA_readData[192]), .A2(n26), .B1(gYMA_readData[208]), 
        .B2(n27), .ZN(n123) );
  AOI22_X2 U17 ( .A1(gYMA_readData[67]), .A2(n14), .B1(gYMA_readData[83]), 
        .B2(n15), .ZN(n83) );
  AOI22_X2 U18 ( .A1(gYMA_readData[66]), .A2(n14), .B1(gYMA_readData[82]), 
        .B2(n15), .ZN(n93) );
  AOI22_X2 U20 ( .A1(gYMA_readData[194]), .A2(n26), .B1(gYMA_readData[210]), 
        .B2(n27), .ZN(n97) );
  AOI22_X2 U21 ( .A1(gYMA_readData[65]), .A2(n14), .B1(gYMA_readData[81]), 
        .B2(n15), .ZN(n103) );
  AOI22_X2 U22 ( .A1(gYMA_readData[193]), .A2(n26), .B1(gYMA_readData[209]), 
        .B2(n27), .ZN(n107) );
  AOI22_X2 U23 ( .A1(gYMA_readData[96]), .A2(n16), .B1(gYMA_readData[112]), 
        .B2(n17), .ZN(n112) );
  AOI22_X2 U24 ( .A1(gYMA_readData[99]), .A2(n16), .B1(gYMA_readData[115]), 
        .B2(n17), .ZN(n82) );
  AOI22_X2 U26 ( .A1(gYMA_readData[98]), .A2(n16), .B1(gYMA_readData[114]), 
        .B2(n17), .ZN(n92) );
  AOI22_X2 U27 ( .A1(gYMA_readData[97]), .A2(n16), .B1(gYMA_readData[113]), 
        .B2(n17), .ZN(n102) );
  AOI22_X2 U28 ( .A1(gYMA_readData[0]), .A2(n10), .B1(gYMA_readData[16]), .B2(
        n11), .ZN(n115) );
  AOI22_X2 U29 ( .A1(gYMA_readData[128]), .A2(n22), .B1(gYMA_readData[144]), 
        .B2(n23), .ZN(n125) );
  AOI22_X2 U31 ( .A1(gYMA_readData[3]), .A2(n10), .B1(gYMA_readData[19]), .B2(
        n11), .ZN(n85) );
  AOI22_X2 U32 ( .A1(gYMA_readData[131]), .A2(n22), .B1(gYMA_readData[147]), 
        .B2(n23), .ZN(n89) );
  AOI22_X2 U33 ( .A1(gYMA_readData[2]), .A2(n10), .B1(gYMA_readData[18]), .B2(
        n11), .ZN(n95) );
  AOI22_X2 U34 ( .A1(gYMA_readData[130]), .A2(n22), .B1(gYMA_readData[146]), 
        .B2(n23), .ZN(n99) );
  AOI22_X2 U35 ( .A1(gYMA_readData[1]), .A2(n10), .B1(gYMA_readData[17]), .B2(
        n11), .ZN(n105) );
  AOI22_X2 U37 ( .A1(gYMA_readData[129]), .A2(n22), .B1(gYMA_readData[145]), 
        .B2(n23), .ZN(n109) );
  AOI22_X2 U38 ( .A1(gYMA_readData[32]), .A2(n12), .B1(gYMA_readData[48]), 
        .B2(n13), .ZN(n114) );
  AOI22_X2 U39 ( .A1(gYMA_readData[160]), .A2(n24), .B1(gYMA_readData[176]), 
        .B2(n25), .ZN(n124) );
  AOI22_X2 U40 ( .A1(gYMA_readData[35]), .A2(n12), .B1(gYMA_readData[51]), 
        .B2(n13), .ZN(n84) );
  AOI22_X2 U42 ( .A1(gYMA_readData[163]), .A2(n24), .B1(gYMA_readData[179]), 
        .B2(n25), .ZN(n88) );
  AOI22_X2 U43 ( .A1(gYMA_readData[34]), .A2(n12), .B1(gYMA_readData[50]), 
        .B2(n13), .ZN(n94) );
  AOI22_X2 U44 ( .A1(gYMA_readData[162]), .A2(n24), .B1(gYMA_readData[178]), 
        .B2(n25), .ZN(n98) );
  AOI22_X2 U45 ( .A1(gYMA_readData[33]), .A2(n12), .B1(gYMA_readData[49]), 
        .B2(n13), .ZN(n104) );
  AOI22_X2 U46 ( .A1(gYMA_readData[161]), .A2(n24), .B1(gYMA_readData[177]), 
        .B2(n25), .ZN(n108) );
  AOI21_X2 U48 ( .B1(n30), .B2(n31), .A(n1), .ZN(gYMA_row_addr1[8]) );
  AOI22_X2 U49 ( .A1(gYMA_readData[232]), .A2(n28), .B1(gYMA_readData[248]), 
        .B2(n29), .ZN(n36) );
  AOI21_X2 U50 ( .B1(n4), .B2(n5), .A(n1), .ZN(gYMA_row_addr1[9]) );
  AOI22_X2 U51 ( .A1(gYMA_readData[233]), .A2(n28), .B1(gYMA_readData[249]), 
        .B2(n29), .ZN(n18) );
  AOI21_X2 U53 ( .B1(n40), .B2(n41), .A(n1), .ZN(gYMA_row_addr1[7]) );
  AOI22_X2 U54 ( .A1(gYMA_readData[231]), .A2(n28), .B1(gYMA_readData[247]), 
        .B2(n29), .ZN(n46) );
  AOI21_X2 U55 ( .B1(n50), .B2(n51), .A(n1), .ZN(gYMA_row_addr1[6]) );
  AOI22_X2 U56 ( .A1(gYMA_readData[230]), .A2(n28), .B1(gYMA_readData[246]), 
        .B2(n29), .ZN(n56) );
  AOI21_X2 U57 ( .B1(n60), .B2(n61), .A(n1), .ZN(gYMA_row_addr1[5]) );
  AOI22_X2 U59 ( .A1(gYMA_readData[229]), .A2(n28), .B1(gYMA_readData[245]), 
        .B2(n29), .ZN(n66) );
  AOI21_X2 U60 ( .B1(n70), .B2(n71), .A(n1), .ZN(gYMA_row_addr1[4]) );
  AOI22_X2 U61 ( .A1(gYMA_readData[228]), .A2(n28), .B1(gYMA_readData[244]), 
        .B2(n29), .ZN(n76) );
  AOI22_X2 U62 ( .A1(gYMA_readData[72]), .A2(n14), .B1(gYMA_readData[88]), 
        .B2(n15), .ZN(n33) );
  AOI22_X2 U64 ( .A1(gYMA_readData[200]), .A2(n26), .B1(gYMA_readData[216]), 
        .B2(n27), .ZN(n37) );
  AOI22_X2 U65 ( .A1(gYMA_readData[73]), .A2(n14), .B1(gYMA_readData[89]), 
        .B2(n15), .ZN(n7) );
  AOI22_X2 U66 ( .A1(gYMA_readData[201]), .A2(n26), .B1(gYMA_readData[217]), 
        .B2(n27), .ZN(n19) );
  AOI22_X2 U67 ( .A1(gYMA_readData[71]), .A2(n14), .B1(gYMA_readData[87]), 
        .B2(n15), .ZN(n43) );
  AOI22_X2 U68 ( .A1(gYMA_readData[199]), .A2(n26), .B1(gYMA_readData[215]), 
        .B2(n27), .ZN(n47) );
  AOI22_X2 U70 ( .A1(gYMA_readData[70]), .A2(n14), .B1(gYMA_readData[86]), 
        .B2(n15), .ZN(n53) );
  AOI22_X2 U71 ( .A1(gYMA_readData[198]), .A2(n26), .B1(gYMA_readData[214]), 
        .B2(n27), .ZN(n57) );
  AOI22_X2 U72 ( .A1(gYMA_readData[69]), .A2(n14), .B1(gYMA_readData[85]), 
        .B2(n15), .ZN(n63) );
  AOI22_X2 U73 ( .A1(gYMA_readData[197]), .A2(n26), .B1(gYMA_readData[213]), 
        .B2(n27), .ZN(n67) );
  AOI22_X2 U75 ( .A1(gYMA_readData[68]), .A2(n14), .B1(gYMA_readData[84]), 
        .B2(n15), .ZN(n73) );
  AOI22_X2 U76 ( .A1(gYMA_readData[196]), .A2(n26), .B1(gYMA_readData[212]), 
        .B2(n27), .ZN(n77) );
  AOI22_X2 U77 ( .A1(gYMA_readData[195]), .A2(n26), .B1(gYMA_readData[211]), 
        .B2(n27), .ZN(n87) );
  AOI22_X2 U78 ( .A1(gYMA_readData[104]), .A2(n16), .B1(gYMA_readData[120]), 
        .B2(n17), .ZN(n32) );
  AOI22_X2 U79 ( .A1(gYMA_readData[105]), .A2(n16), .B1(gYMA_readData[121]), 
        .B2(n17), .ZN(n6) );
  AOI22_X2 U81 ( .A1(gYMA_readData[103]), .A2(n16), .B1(gYMA_readData[119]), 
        .B2(n17), .ZN(n42) );
  AOI22_X2 U82 ( .A1(gYMA_readData[102]), .A2(n16), .B1(gYMA_readData[118]), 
        .B2(n17), .ZN(n52) );
  AOI22_X2 U83 ( .A1(gYMA_readData[101]), .A2(n16), .B1(gYMA_readData[117]), 
        .B2(n17), .ZN(n62) );
  AOI22_X2 U84 ( .A1(gYMA_readData[100]), .A2(n16), .B1(gYMA_readData[116]), 
        .B2(n17), .ZN(n72) );
  AOI22_X2 U86 ( .A1(gYMA_readData[8]), .A2(n10), .B1(gYMA_readData[24]), .B2(
        n11), .ZN(n35) );
  AOI22_X2 U87 ( .A1(gYMA_readData[136]), .A2(n22), .B1(gYMA_readData[152]), 
        .B2(n23), .ZN(n39) );
  AOI22_X2 U88 ( .A1(gYMA_readData[9]), .A2(n10), .B1(gYMA_readData[25]), .B2(
        n11), .ZN(n9) );
  AOI22_X2 U89 ( .A1(gYMA_readData[137]), .A2(n22), .B1(gYMA_readData[153]), 
        .B2(n23), .ZN(n21) );
  AOI22_X2 U90 ( .A1(gYMA_readData[7]), .A2(n10), .B1(gYMA_readData[23]), .B2(
        n11), .ZN(n45) );
  AOI22_X2 U92 ( .A1(gYMA_readData[135]), .A2(n22), .B1(gYMA_readData[151]), 
        .B2(n23), .ZN(n49) );
  AOI22_X2 U93 ( .A1(gYMA_readData[6]), .A2(n10), .B1(gYMA_readData[22]), .B2(
        n11), .ZN(n55) );
  AOI22_X2 U94 ( .A1(gYMA_readData[134]), .A2(n22), .B1(gYMA_readData[150]), 
        .B2(n23), .ZN(n59) );
  AOI22_X2 U95 ( .A1(gYMA_readData[5]), .A2(n10), .B1(gYMA_readData[21]), .B2(
        n11), .ZN(n65) );
  AOI22_X2 U97 ( .A1(gYMA_readData[133]), .A2(n22), .B1(gYMA_readData[149]), 
        .B2(n23), .ZN(n69) );
  AOI22_X2 U98 ( .A1(gYMA_readData[4]), .A2(n10), .B1(gYMA_readData[20]), .B2(
        n11), .ZN(n75) );
  AOI22_X2 U99 ( .A1(gYMA_readData[132]), .A2(n22), .B1(gYMA_readData[148]), 
        .B2(n23), .ZN(n79) );
  AOI22_X2 U100 ( .A1(gYMA_readData[40]), .A2(n12), .B1(gYMA_readData[56]), 
        .B2(n13), .ZN(n34) );
  AOI22_X2 U101 ( .A1(gYMA_readData[168]), .A2(n24), .B1(gYMA_readData[184]), 
        .B2(n25), .ZN(n38) );
  AOI22_X2 U103 ( .A1(gYMA_readData[41]), .A2(n12), .B1(gYMA_readData[57]), 
        .B2(n13), .ZN(n8) );
  AOI22_X2 U104 ( .A1(gYMA_readData[169]), .A2(n24), .B1(gYMA_readData[185]), 
        .B2(n25), .ZN(n20) );
  AOI22_X2 U105 ( .A1(gYMA_readData[39]), .A2(n12), .B1(gYMA_readData[55]), 
        .B2(n13), .ZN(n44) );
  AOI22_X2 U106 ( .A1(gYMA_readData[167]), .A2(n24), .B1(gYMA_readData[183]), 
        .B2(n25), .ZN(n48) );
  AOI22_X2 U108 ( .A1(gYMA_readData[38]), .A2(n12), .B1(gYMA_readData[54]), 
        .B2(n13), .ZN(n54) );
  AOI22_X2 U109 ( .A1(gYMA_readData[166]), .A2(n24), .B1(gYMA_readData[182]), 
        .B2(n25), .ZN(n58) );
  AOI22_X2 U110 ( .A1(gYMA_readData[37]), .A2(n12), .B1(gYMA_readData[53]), 
        .B2(n13), .ZN(n64) );
  AOI22_X2 U112 ( .A1(gYMA_readData[165]), .A2(n24), .B1(gYMA_readData[181]), 
        .B2(n25), .ZN(n68) );
  AOI22_X2 U116 ( .A1(gYMA_readData[36]), .A2(n12), .B1(gYMA_readData[52]), 
        .B2(n13), .ZN(n74) );
  AOI22_X2 U119 ( .A1(gYMA_readData[164]), .A2(n24), .B1(gYMA_readData[180]), 
        .B2(n25), .ZN(n78) );
  INV_X4 U120 ( .A(readEnable), .ZN(n1) );
  AND2_X4 U121 ( .A1(n127), .A2(n121), .ZN(n28) );
  AND2_X4 U122 ( .A1(n126), .A2(n121), .ZN(n29) );
  AND2_X4 U123 ( .A1(n127), .A2(n120), .ZN(n26) );
  AND2_X4 U124 ( .A1(n126), .A2(n120), .ZN(n27) );
  AND2_X4 U125 ( .A1(n127), .A2(n119), .ZN(n24) );
  AND2_X4 U127 ( .A1(n126), .A2(n119), .ZN(n25) );
  AND2_X4 U129 ( .A1(n127), .A2(n117), .ZN(n22) );
  AND2_X4 U130 ( .A1(n126), .A2(n117), .ZN(n23) );
  AND2_X4 U132 ( .A1(n121), .A2(n118), .ZN(n16) );
  AND2_X4 U133 ( .A1(n121), .A2(n116), .ZN(n17) );
  AND2_X4 U135 ( .A1(n120), .A2(n118), .ZN(n14) );
  AND2_X4 U136 ( .A1(n120), .A2(n116), .ZN(n15) );
  AND2_X4 U137 ( .A1(n119), .A2(n118), .ZN(n12) );
  AND2_X4 U138 ( .A1(n119), .A2(n116), .ZN(n13) );
  AND2_X4 U139 ( .A1(n117), .A2(n118), .ZN(n10) );
  AND2_X4 U140 ( .A1(n116), .A2(n117), .ZN(n11) );
endmodule


module yAddrDecodr ( clock, reset, yAD_enable, yAD_readRowNum, yAD_readRowData, 
        yAD_outAddr1, yAD_outAddr2, yAD_dataOutNextCycle );
  input [15:0] yAD_readRowNum;
  input [255:0] yAD_readRowData;
  output [10:0] yAD_outAddr1;
  output [10:0] yAD_outAddr2;
  input clock, reset, yAD_enable;
  output yAD_dataOutNextCycle;
  wire   n54, n116, n118, U3_U1_DATA2_0, U3_U1_DATA2_1, U3_U1_DATA2_2,
         U3_U1_DATA2_3, U3_U1_DATA2_4, U3_U1_DATA2_5, U3_U1_DATA2_6,
         U3_U1_DATA2_7, U3_U1_DATA2_8, U3_U1_DATA2_9, U3_U2_Z_0, U5_Z_0,
         U5_Z_1, U5_Z_2, U5_Z_3, U5_Z_4, U5_Z_5, U5_Z_6, U5_Z_7, U5_Z_8,
         U5_Z_9, U5_Z_10, U5_DATA2_2, U5_DATA2_3, U5_DATA2_4, U5_DATA2_5,
         U5_DATA2_6, U5_DATA2_7, U5_DATA2_8, U5_DATA2_9, U5_DATA2_10, U4_Z_0,
         U4_Z_1, U4_Z_2, U4_Z_3, U4_Z_4, U4_Z_5, U4_Z_6, U4_Z_7, U4_Z_8,
         U4_Z_9, U4_Z_10, U4_DATA3_0, U4_DATA3_1, U4_DATA3_2, U4_DATA3_3,
         U4_DATA3_4, U4_DATA3_5, U4_DATA3_6, U4_DATA3_7, U4_DATA3_8,
         U4_DATA3_9, U4_DATA3_10, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n13, n14, n16, n17, n18, n19, n20, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n43, n44,
         n46, n47, n48, n49, n50, n51, n52, n53, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n90, n91, n92, n93, n94, n95, n96, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, SYNOPSYS_UNCONNECTED_1;
  wire   [115:100] n;
  wire   [9:2] r313_carry;
  wire   [9:3] add_52_carry;

  getYMatAddress gY2 ( .readEnable(n116), .gYMA_row(n), .gYMA_readData(
        yAD_readRowData), .gYMA_row_addr1({SYNOPSYS_UNCONNECTED_1, 
        U3_U1_DATA2_9, U3_U1_DATA2_8, U3_U1_DATA2_7, U3_U1_DATA2_6, 
        U3_U1_DATA2_5, U3_U1_DATA2_4, U3_U1_DATA2_3, U3_U1_DATA2_2, 
        U3_U1_DATA2_1, U3_U1_DATA2_0}) );
  FA_X1 r313_U1_1 ( .A(n31), .B(n455), .CI(n435), .CO(r313_carry[2]), .S(
        U4_DATA3_1) );
  DFF_X1 temp_bit_reg ( .D(n54), .CK(clock), .Q(n118) );
  DFF_X1 reg_readEn_reg ( .D(n43), .CK(clock), .Q(n116) );
  DFF_X1 yAD_dataOutNextCycle_reg ( .D(n456), .CK(clock), .Q(
        yAD_dataOutNextCycle) );
  DFF_X1 temp_oldRow_reg_15_ ( .D(n2), .CK(clock), .Q(n[115]) );
  DFF_X1 temp_oldRow_reg_14_ ( .D(n3), .CK(clock), .Q(n[114]) );
  DFF_X1 temp_oldRow_reg_13_ ( .D(n4), .CK(clock), .Q(n[113]) );
  DFF_X1 temp_oldRow_reg_12_ ( .D(n5), .CK(clock), .Q(n[112]) );
  DFF_X1 temp_oldRow_reg_11_ ( .D(n6), .CK(clock), .Q(n[111]) );
  DFF_X1 temp_oldRow_reg_10_ ( .D(n7), .CK(clock), .Q(n[110]) );
  DFF_X1 temp_oldRow_reg_9_ ( .D(n8), .CK(clock), .Q(n[109]) );
  DFF_X1 temp_oldRow_reg_8_ ( .D(n9), .CK(clock), .Q(n[108]) );
  DFF_X1 temp_oldRow_reg_7_ ( .D(n10), .CK(clock), .Q(n[107]) );
  DFF_X1 temp_oldRow_reg_6_ ( .D(n11), .CK(clock), .Q(n[106]) );
  DFF_X1 temp_oldRow_reg_5_ ( .D(n13), .CK(clock), .Q(n[105]) );
  DFF_X1 temp_oldRow_reg_4_ ( .D(n14), .CK(clock), .Q(n[104]) );
  DFF_X1 temp_oldRow_reg_3_ ( .D(n16), .CK(clock), .Q(n[103]) );
  DFF_X1 temp_oldRow_reg_2_ ( .D(n17), .CK(clock), .Q(n[102]) );
  DFF_X1 temp_oldRow_reg_1_ ( .D(n18), .CK(clock), .Q(n[101]) );
  DFF_X1 temp_oldRow_reg_0_ ( .D(n19), .CK(clock), .Q(n[100]) );
  DFF_X1 yAD_outAddr1_reg_1_ ( .D(U5_Z_1), .CK(clock), .Q(yAD_outAddr1[1]), 
        .QN(n437) );
  DFF_X1 yAD_outAddr1_reg_2_ ( .D(U5_Z_2), .CK(clock), .Q(yAD_outAddr1[2]) );
  DFF_X1 yAD_outAddr1_reg_3_ ( .D(U5_Z_3), .CK(clock), .Q(yAD_outAddr1[3]) );
  DFF_X1 yAD_outAddr1_reg_4_ ( .D(U5_Z_4), .CK(clock), .Q(yAD_outAddr1[4]) );
  DFF_X1 yAD_outAddr1_reg_5_ ( .D(U5_Z_5), .CK(clock), .Q(yAD_outAddr1[5]) );
  DFF_X1 yAD_outAddr1_reg_6_ ( .D(U5_Z_6), .CK(clock), .Q(yAD_outAddr1[6]) );
  DFF_X1 yAD_outAddr1_reg_7_ ( .D(U5_Z_7), .CK(clock), .Q(yAD_outAddr1[7]) );
  DFF_X1 yAD_outAddr1_reg_8_ ( .D(U5_Z_8), .CK(clock), .Q(yAD_outAddr1[8]) );
  DFF_X1 yAD_outAddr1_reg_9_ ( .D(U5_Z_9), .CK(clock), .Q(yAD_outAddr1[9]) );
  DFF_X1 yAD_outAddr1_reg_10_ ( .D(U5_Z_10), .CK(clock), .Q(yAD_outAddr1[10])
         );
  DFF_X1 yAD_outAddr1_reg_0_ ( .D(U5_Z_0), .CK(clock), .Q(yAD_outAddr1[0]) );
  DFF_X1 yAD_outAddr2_reg_0_ ( .D(U4_Z_0), .CK(clock), .Q(yAD_outAddr2[0]) );
  DFF_X1 yAD_outAddr2_reg_1_ ( .D(U4_Z_1), .CK(clock), .Q(yAD_outAddr2[1]) );
  DFF_X1 yAD_outAddr2_reg_2_ ( .D(U4_Z_2), .CK(clock), .Q(yAD_outAddr2[2]) );
  DFF_X1 yAD_outAddr2_reg_3_ ( .D(U4_Z_3), .CK(clock), .Q(yAD_outAddr2[3]) );
  DFF_X1 yAD_outAddr2_reg_4_ ( .D(U4_Z_4), .CK(clock), .Q(yAD_outAddr2[4]) );
  DFF_X1 yAD_outAddr2_reg_5_ ( .D(U4_Z_5), .CK(clock), .Q(yAD_outAddr2[5]) );
  DFF_X1 yAD_outAddr2_reg_6_ ( .D(U4_Z_6), .CK(clock), .Q(yAD_outAddr2[6]) );
  DFF_X1 yAD_outAddr2_reg_7_ ( .D(U4_Z_7), .CK(clock), .Q(yAD_outAddr2[7]) );
  DFF_X1 yAD_outAddr2_reg_8_ ( .D(U4_Z_8), .CK(clock), .Q(yAD_outAddr2[8]) );
  DFF_X1 yAD_outAddr2_reg_9_ ( .D(U4_Z_9), .CK(clock), .Q(yAD_outAddr2[9]) );
  DFF_X1 yAD_outAddr2_reg_10_ ( .D(U4_Z_10), .CK(clock), .Q(yAD_outAddr2[10])
         );
  AOI221_X2 U3 ( .B1(yAD_readRowNum[0]), .B2(n456), .C1(n20), .C2(n[100]), .A(
        n48), .ZN(n47) );
  AOI221_X2 U4 ( .B1(yAD_readRowNum[1]), .B2(n456), .C1(n20), .C2(n[101]), .A(
        n48), .ZN(n49) );
  AOI221_X2 U5 ( .B1(yAD_readRowNum[2]), .B2(n456), .C1(n20), .C2(n[102]), .A(
        n48), .ZN(n50) );
  AOI221_X2 U8 ( .B1(yAD_readRowNum[3]), .B2(n456), .C1(n20), .C2(n[103]), .A(
        n48), .ZN(n51) );
  AOI221_X2 U9 ( .B1(yAD_readRowNum[4]), .B2(n456), .C1(n20), .C2(n[104]), .A(
        n48), .ZN(n52) );
  AOI221_X2 U10 ( .B1(yAD_readRowNum[5]), .B2(n456), .C1(n20), .C2(n[105]), 
        .A(n48), .ZN(n53) );
  AOI221_X2 U11 ( .B1(yAD_readRowNum[6]), .B2(n456), .C1(n20), .C2(n[106]), 
        .A(n48), .ZN(n55) );
  AOI221_X2 U12 ( .B1(yAD_readRowNum[7]), .B2(n456), .C1(n20), .C2(n[107]), 
        .A(n48), .ZN(n56) );
  AOI221_X2 U13 ( .B1(yAD_readRowNum[8]), .B2(n456), .C1(n20), .C2(n[108]), 
        .A(n48), .ZN(n57) );
  AOI221_X2 U14 ( .B1(yAD_readRowNum[9]), .B2(n456), .C1(n20), .C2(n[109]), 
        .A(n48), .ZN(n58) );
  AOI221_X2 U15 ( .B1(yAD_readRowNum[10]), .B2(n456), .C1(n20), .C2(n[110]), 
        .A(n48), .ZN(n59) );
  NAND2_X2 U21 ( .A1(n66), .A2(n43), .ZN(n54) );
  NOR2_X2 U22 ( .A1(n68), .A2(n69), .ZN(n66) );
  OAI221_X2 U41 ( .B1(yAD_outAddr1[1]), .B2(n44), .C1(n46), .C2(n67), .A(n79), 
        .ZN(U5_Z_1) );
  NOR3_X2 U46 ( .A1(n455), .A2(n118), .A3(n48), .ZN(n69) );
  NAND2_X2 U47 ( .A1(n43), .A2(n67), .ZN(n65) );
  NAND3_X2 U48 ( .A1(n43), .A2(U3_U2_Z_0), .A3(n118), .ZN(n67) );
  AND3_X2 U62 ( .A1(n96), .A2(yAD_readRowNum[10]), .A3(yAD_readRowNum[11]), 
        .ZN(n95) );
  AND3_X2 U63 ( .A1(yAD_readRowNum[0]), .A2(yAD_enable), .A3(yAD_readRowNum[1]), .ZN(n96) );
  AND4_X2 U64 ( .A1(yAD_readRowNum[12]), .A2(yAD_readRowNum[13]), .A3(
        yAD_readRowNum[14]), .A4(yAD_readRowNum[15]), .ZN(n94) );
  AND4_X2 U65 ( .A1(yAD_readRowNum[2]), .A2(yAD_readRowNum[3]), .A3(
        yAD_readRowNum[4]), .A4(yAD_readRowNum[5]), .ZN(n93) );
  AND4_X2 U66 ( .A1(yAD_readRowNum[6]), .A2(yAD_readRowNum[7]), .A3(
        yAD_readRowNum[8]), .A4(yAD_readRowNum[9]), .ZN(n92) );
  INV_X4 U67 ( .A(n69), .ZN(n1) );
  INV_X4 U68 ( .A(n64), .ZN(n2) );
  INV_X4 U69 ( .A(n63), .ZN(n3) );
  INV_X4 U70 ( .A(n62), .ZN(n4) );
  INV_X4 U71 ( .A(n61), .ZN(n5) );
  INV_X4 U72 ( .A(n60), .ZN(n6) );
  INV_X4 U73 ( .A(n59), .ZN(n7) );
  INV_X4 U74 ( .A(n58), .ZN(n8) );
  INV_X4 U75 ( .A(n57), .ZN(n9) );
  INV_X4 U76 ( .A(n56), .ZN(n10) );
  INV_X4 U77 ( .A(n55), .ZN(n11) );
  INV_X4 U78 ( .A(n53), .ZN(n13) );
  INV_X4 U79 ( .A(n52), .ZN(n14) );
  INV_X4 U80 ( .A(n51), .ZN(n16) );
  INV_X4 U81 ( .A(n50), .ZN(n17) );
  INV_X4 U82 ( .A(n49), .ZN(n18) );
  INV_X4 U83 ( .A(n47), .ZN(n19) );
  INV_X4 U87 ( .A(n81), .ZN(n23) );
  INV_X4 U88 ( .A(n82), .ZN(n24) );
  INV_X4 U89 ( .A(n83), .ZN(n25) );
  INV_X4 U90 ( .A(n84), .ZN(n26) );
  INV_X4 U91 ( .A(n85), .ZN(n27) );
  INV_X4 U92 ( .A(n86), .ZN(n28) );
  INV_X4 U93 ( .A(n87), .ZN(n29) );
  INV_X4 U94 ( .A(n88), .ZN(n30) );
  INV_X4 U95 ( .A(n90), .ZN(n31) );
  INV_X4 U96 ( .A(n91), .ZN(n32) );
  INV_X4 U97 ( .A(U3_U1_DATA2_0), .ZN(n33) );
  INV_X4 U98 ( .A(U3_U1_DATA2_2), .ZN(n34) );
  INV_X4 U99 ( .A(U3_U1_DATA2_3), .ZN(n35) );
  INV_X4 U100 ( .A(U3_U1_DATA2_4), .ZN(n36) );
  INV_X4 U101 ( .A(U3_U1_DATA2_5), .ZN(n37) );
  INV_X4 U102 ( .A(U3_U1_DATA2_6), .ZN(n38) );
  INV_X4 U103 ( .A(U3_U1_DATA2_7), .ZN(n39) );
  INV_X4 U104 ( .A(U3_U1_DATA2_8), .ZN(n40) );
  INV_X4 U105 ( .A(U3_U1_DATA2_9), .ZN(n41) );
  INV_X4 U108 ( .A(n68), .ZN(n44) );
  INV_X4 U110 ( .A(yAD_readRowNum[5]), .ZN(n46) );
  OR2_X1 U111 ( .A1(U4_DATA3_9), .A2(n65), .ZN(U4_Z_9) );
  OR2_X1 U112 ( .A1(U4_DATA3_8), .A2(n65), .ZN(U4_Z_8) );
  OR2_X1 U113 ( .A1(U4_DATA3_7), .A2(n65), .ZN(U4_Z_7) );
  OR2_X1 U114 ( .A1(U4_DATA3_6), .A2(n65), .ZN(U4_Z_6) );
  OR2_X1 U115 ( .A1(U4_DATA3_5), .A2(n65), .ZN(U4_Z_5) );
  OR2_X1 U116 ( .A1(U4_DATA3_4), .A2(n65), .ZN(U4_Z_4) );
  OR2_X1 U117 ( .A1(U4_DATA3_3), .A2(n65), .ZN(U4_Z_3) );
  OR2_X1 U118 ( .A1(U4_DATA3_2), .A2(n65), .ZN(U4_Z_2) );
  OR2_X1 U119 ( .A1(U4_DATA3_10), .A2(n65), .ZN(U4_Z_10) );
  OR2_X1 U120 ( .A1(U4_DATA3_1), .A2(n65), .ZN(U4_Z_1) );
  OR2_X1 U121 ( .A1(U4_DATA3_0), .A2(n65), .ZN(U4_Z_0) );
  AND2_X4 U6 ( .A1(U3_U2_Z_0), .A2(n32), .ZN(n435) );
  AND2_X4 U7 ( .A1(n455), .A2(yAD_outAddr2[10]), .ZN(n436) );
  INV_X4 U16 ( .A(n65), .ZN(n20) );
  INV_X4 U17 ( .A(n67), .ZN(n456) );
  NOR2_X2 U18 ( .A1(n48), .A2(U3_U2_Z_0), .ZN(n68) );
  INV_X4 U19 ( .A(n48), .ZN(n43) );
  AOI22_X2 U20 ( .A1(n455), .A2(yAD_outAddr2[1]), .B1(U3_U2_Z_0), .B2(
        U3_U1_DATA2_1), .ZN(n90) );
  INV_X4 U23 ( .A(U3_U2_Z_0), .ZN(n455) );
  NAND4_X2 U24 ( .A1(n92), .A2(n93), .A3(n94), .A4(n95), .ZN(U3_U2_Z_0) );
  AOI22_X2 U25 ( .A1(n455), .A2(yAD_outAddr2[3]), .B1(U3_U2_Z_0), .B2(
        U3_U1_DATA2_3), .ZN(n87) );
  AOI22_X2 U26 ( .A1(n455), .A2(yAD_outAddr2[0]), .B1(U3_U2_Z_0), .B2(
        U3_U1_DATA2_0), .ZN(n91) );
  AOI22_X2 U27 ( .A1(n455), .A2(yAD_outAddr2[2]), .B1(U3_U2_Z_0), .B2(
        U3_U1_DATA2_2), .ZN(n88) );
  AOI22_X2 U28 ( .A1(n455), .A2(yAD_outAddr2[5]), .B1(U3_U2_Z_0), .B2(
        U3_U1_DATA2_5), .ZN(n85) );
  AOI22_X2 U29 ( .A1(n455), .A2(yAD_outAddr2[7]), .B1(U3_U2_Z_0), .B2(
        U3_U1_DATA2_7), .ZN(n83) );
  AOI22_X2 U30 ( .A1(n455), .A2(yAD_outAddr2[8]), .B1(U3_U2_Z_0), .B2(
        U3_U1_DATA2_8), .ZN(n82) );
  AOI22_X2 U31 ( .A1(n455), .A2(yAD_outAddr2[9]), .B1(U3_U2_Z_0), .B2(
        U3_U1_DATA2_9), .ZN(n81) );
  AOI22_X2 U32 ( .A1(n455), .A2(yAD_outAddr2[4]), .B1(U3_U2_Z_0), .B2(
        U3_U1_DATA2_4), .ZN(n86) );
  AOI22_X2 U33 ( .A1(n455), .A2(yAD_outAddr2[6]), .B1(U3_U2_Z_0), .B2(
        U3_U1_DATA2_6), .ZN(n84) );
  NAND2_X2 U34 ( .A1(reset), .A2(yAD_enable), .ZN(n48) );
  AOI22_X2 U35 ( .A1(U5_DATA2_10), .A2(n68), .B1(n456), .B2(yAD_readRowNum[14]), .ZN(n78) );
  OAI211_X2 U36 ( .C1(n1), .C2(n41), .A(n43), .B(n70), .ZN(U5_Z_9) );
  AOI22_X2 U37 ( .A1(U5_DATA2_9), .A2(n68), .B1(n456), .B2(yAD_readRowNum[13]), 
        .ZN(n70) );
  OAI211_X2 U38 ( .C1(n1), .C2(n40), .A(n43), .B(n71), .ZN(U5_Z_8) );
  AOI22_X2 U39 ( .A1(U5_DATA2_8), .A2(n68), .B1(n456), .B2(yAD_readRowNum[12]), 
        .ZN(n71) );
  OAI211_X2 U40 ( .C1(n1), .C2(n39), .A(n43), .B(n72), .ZN(U5_Z_7) );
  AOI22_X2 U42 ( .A1(U5_DATA2_7), .A2(n68), .B1(n456), .B2(yAD_readRowNum[11]), 
        .ZN(n72) );
  OAI211_X2 U43 ( .C1(n1), .C2(n38), .A(n43), .B(n73), .ZN(U5_Z_6) );
  AOI22_X2 U44 ( .A1(U5_DATA2_6), .A2(n68), .B1(n456), .B2(yAD_readRowNum[10]), 
        .ZN(n73) );
  OAI211_X2 U45 ( .C1(n1), .C2(n37), .A(n43), .B(n74), .ZN(U5_Z_5) );
  AOI22_X2 U49 ( .A1(U5_DATA2_5), .A2(n68), .B1(n456), .B2(yAD_readRowNum[9]), 
        .ZN(n74) );
  OAI211_X2 U50 ( .C1(n1), .C2(n36), .A(n43), .B(n75), .ZN(U5_Z_4) );
  AOI22_X2 U51 ( .A1(U5_DATA2_4), .A2(n68), .B1(n456), .B2(yAD_readRowNum[8]), 
        .ZN(n75) );
  OAI211_X2 U52 ( .C1(n1), .C2(n35), .A(n43), .B(n76), .ZN(U5_Z_3) );
  AOI22_X2 U53 ( .A1(U5_DATA2_3), .A2(n68), .B1(n456), .B2(yAD_readRowNum[7]), 
        .ZN(n76) );
  OAI211_X2 U54 ( .C1(n1), .C2(n34), .A(n43), .B(n77), .ZN(U5_Z_2) );
  AOI22_X2 U55 ( .A1(U5_DATA2_2), .A2(n68), .B1(n456), .B2(yAD_readRowNum[6]), 
        .ZN(n77) );
  OAI211_X2 U56 ( .C1(n1), .C2(n33), .A(n43), .B(n80), .ZN(U5_Z_0) );
  AOI22_X2 U57 ( .A1(yAD_outAddr1[0]), .A2(n68), .B1(n456), .B2(
        yAD_readRowNum[4]), .ZN(n80) );
  AOI21_X2 U58 ( .B1(U3_U1_DATA2_1), .B2(n69), .A(n48), .ZN(n79) );
  AOI22_X2 U59 ( .A1(n20), .A2(n[111]), .B1(yAD_readRowNum[11]), .B2(n456), 
        .ZN(n60) );
  AOI22_X2 U60 ( .A1(n20), .A2(n[112]), .B1(yAD_readRowNum[12]), .B2(n456), 
        .ZN(n61) );
  AOI22_X2 U61 ( .A1(n20), .A2(n[113]), .B1(yAD_readRowNum[13]), .B2(n456), 
        .ZN(n62) );
  AOI22_X2 U84 ( .A1(n20), .A2(n[114]), .B1(yAD_readRowNum[14]), .B2(n456), 
        .ZN(n63) );
  AOI22_X2 U85 ( .A1(n20), .A2(n[115]), .B1(yAD_readRowNum[15]), .B2(n456), 
        .ZN(n64) );
  XNOR2_X2 U86 ( .A(U3_U2_Z_0), .B(n91), .ZN(U4_DATA3_0) );
  INV_X4 U106 ( .A(r313_carry[2]), .ZN(n438) );
  XNOR2_X2 U107 ( .A(n30), .B(n438), .ZN(U4_DATA3_2) );
  NAND2_X2 U109 ( .A1(n30), .A2(r313_carry[2]), .ZN(n439) );
  INV_X4 U122 ( .A(n439), .ZN(r313_carry[3]) );
  XNOR2_X2 U123 ( .A(n29), .B(n439), .ZN(U4_DATA3_3) );
  NAND2_X2 U124 ( .A1(n29), .A2(r313_carry[3]), .ZN(n440) );
  INV_X4 U125 ( .A(n440), .ZN(r313_carry[4]) );
  XNOR2_X2 U126 ( .A(n28), .B(n440), .ZN(U4_DATA3_4) );
  NAND2_X2 U127 ( .A1(n28), .A2(r313_carry[4]), .ZN(n441) );
  INV_X4 U128 ( .A(n441), .ZN(r313_carry[5]) );
  XNOR2_X2 U129 ( .A(n27), .B(n441), .ZN(U4_DATA3_5) );
  NAND2_X2 U130 ( .A1(n27), .A2(r313_carry[5]), .ZN(n442) );
  INV_X4 U131 ( .A(n442), .ZN(r313_carry[6]) );
  XNOR2_X2 U132 ( .A(n26), .B(n442), .ZN(U4_DATA3_6) );
  NAND2_X2 U133 ( .A1(n26), .A2(r313_carry[6]), .ZN(n443) );
  INV_X4 U134 ( .A(n443), .ZN(r313_carry[7]) );
  XNOR2_X2 U135 ( .A(n25), .B(n443), .ZN(U4_DATA3_7) );
  NAND2_X2 U136 ( .A1(n25), .A2(r313_carry[7]), .ZN(n444) );
  INV_X4 U137 ( .A(n444), .ZN(r313_carry[8]) );
  XNOR2_X2 U138 ( .A(n24), .B(n444), .ZN(U4_DATA3_8) );
  NAND2_X2 U139 ( .A1(n24), .A2(r313_carry[8]), .ZN(n445) );
  INV_X4 U140 ( .A(n445), .ZN(r313_carry[9]) );
  XNOR2_X2 U141 ( .A(n23), .B(n445), .ZN(U4_DATA3_9) );
  NAND2_X2 U142 ( .A1(n23), .A2(r313_carry[9]), .ZN(n446) );
  XNOR2_X2 U143 ( .A(n436), .B(n446), .ZN(U4_DATA3_10) );
  XNOR2_X2 U144 ( .A(yAD_outAddr1[2]), .B(n437), .ZN(U5_DATA2_2) );
  NAND2_X2 U145 ( .A1(yAD_outAddr1[2]), .A2(yAD_outAddr1[1]), .ZN(n447) );
  INV_X4 U146 ( .A(n447), .ZN(add_52_carry[3]) );
  XNOR2_X2 U147 ( .A(yAD_outAddr1[3]), .B(n447), .ZN(U5_DATA2_3) );
  NAND2_X2 U148 ( .A1(yAD_outAddr1[3]), .A2(add_52_carry[3]), .ZN(n448) );
  INV_X4 U149 ( .A(n448), .ZN(add_52_carry[4]) );
  XNOR2_X2 U150 ( .A(yAD_outAddr1[4]), .B(n448), .ZN(U5_DATA2_4) );
  NAND2_X2 U151 ( .A1(yAD_outAddr1[4]), .A2(add_52_carry[4]), .ZN(n449) );
  INV_X4 U152 ( .A(n449), .ZN(add_52_carry[5]) );
  XNOR2_X2 U153 ( .A(yAD_outAddr1[5]), .B(n449), .ZN(U5_DATA2_5) );
  NAND2_X2 U154 ( .A1(yAD_outAddr1[5]), .A2(add_52_carry[5]), .ZN(n450) );
  INV_X4 U155 ( .A(n450), .ZN(add_52_carry[6]) );
  XNOR2_X2 U156 ( .A(yAD_outAddr1[6]), .B(n450), .ZN(U5_DATA2_6) );
  NAND2_X2 U157 ( .A1(yAD_outAddr1[6]), .A2(add_52_carry[6]), .ZN(n451) );
  INV_X4 U158 ( .A(n451), .ZN(add_52_carry[7]) );
  XNOR2_X2 U159 ( .A(yAD_outAddr1[7]), .B(n451), .ZN(U5_DATA2_7) );
  NAND2_X2 U160 ( .A1(yAD_outAddr1[7]), .A2(add_52_carry[7]), .ZN(n452) );
  INV_X4 U161 ( .A(n452), .ZN(add_52_carry[8]) );
  XNOR2_X2 U162 ( .A(yAD_outAddr1[8]), .B(n452), .ZN(U5_DATA2_8) );
  NAND2_X2 U163 ( .A1(yAD_outAddr1[8]), .A2(add_52_carry[8]), .ZN(n453) );
  INV_X4 U164 ( .A(n453), .ZN(add_52_carry[9]) );
  XNOR2_X2 U165 ( .A(yAD_outAddr1[9]), .B(n453), .ZN(U5_DATA2_9) );
  NAND2_X2 U166 ( .A1(yAD_outAddr1[9]), .A2(add_52_carry[9]), .ZN(n454) );
  XNOR2_X2 U167 ( .A(yAD_outAddr1[10]), .B(n454), .ZN(U5_DATA2_10) );
  NAND2_X2 U168 ( .A1(n43), .A2(n78), .ZN(U5_Z_10) );
endmodule


module updateYcomputation ( clock, reset, computationEnable, uYc_chgTxt_row, 
        uYc_chgTxt_col, uYc_chgTxt_real, uYc_chgTxt_img, uYc_ySRAM_rowRead1, 
        uYc_ySRAM_rowRead2, uYc_yMatAddrOut1, uYc_yMatAddrOut2, 
        uYc_dataPathDoneFlag, uYc_filtYopDone, uYc_opYval, uYc_writeDiagAddr, 
        uYc_writeNonDiagAddr, uYc_writeDiagOneHot, uYc_writeNonDiagOneHot, 
        uYC_op_fpIn1, uYC_op_fpIn2, uYC_op_fpMode, uYC_in_fpOut );
  input [15:0] uYc_chgTxt_row;
  input [15:0] uYc_chgTxt_col;
  input [23:0] uYc_chgTxt_real;
  input [23:0] uYc_chgTxt_img;
  input [255:0] uYc_ySRAM_rowRead1;
  input [255:0] uYc_ySRAM_rowRead2;
  output [10:0] uYc_yMatAddrOut1;
  output [10:0] uYc_yMatAddrOut2;
  output [47:0] uYc_opYval;
  output [10:0] uYc_writeDiagAddr;
  output [10:0] uYc_writeNonDiagAddr;
  output [3:0] uYc_writeDiagOneHot;
  output [3:0] uYc_writeNonDiagOneHot;
  output [47:0] uYC_op_fpIn1;
  output [47:0] uYC_op_fpIn2;
  input [47:0] uYC_in_fpOut;
  input clock, reset, computationEnable;
  output uYc_dataPathDoneFlag, uYc_filtYopDone, uYC_op_fpMode;
  wire   wire_execEnable, wire_dataOuNxtCycle, wire_execDoneFlag,
         wire_yAD_Enable;
  wire   [47:0] uYc_filtYval1;
  wire   [47:0] uYc_filtYval2;
  wire   [15:0] uYc_opRowNum_from_filtY;

  updateY_datapath unit_dataPath1 ( .clock(clock), .reset(reset), 
        .executeEnableBit(wire_execEnable), .yInVal1(uYc_filtYval1), .yInVal2(
        uYc_filtYval2), .op_yWriteVal(uYc_opYval), .op_DoneFlag(
        uYc_dataPathDoneFlag), .op_ExDoneFlag(wire_execDoneFlag), 
        .op_CPDoneFlag(uYc_filtYopDone), .op_fpIn1(uYC_op_fpIn1), .op_fpIn2(
        uYC_op_fpIn2), .op_fpMode(uYC_op_fpMode), .in_fpOut(uYC_in_fpOut) );
  updateY_control unit_controlY1 ( .clock(clock), .reset(reset), .exModDone(
        wire_execDoneFlag), .chng_row(uYc_chgTxt_row), .chng_col(
        uYc_chgTxt_col), .chng_real(uYc_chgTxt_real), .chng_img(uYc_chgTxt_img), .dpModDoneFlag(uYc_dataPathDoneFlag), .ymem_data1(uYc_ySRAM_rowRead1), 
        .ymem_data2(uYc_ySRAM_rowRead2), .filt_EN(computationEnable), 
        .yMemDataReadyNextCycle(wire_dataOuNxtCycle), .yAddrIn1(
        uYc_yMatAddrOut1), .yAddrIn2(uYc_yMatAddrOut2), .op_y_row(
        uYc_opRowNum_from_filtY), .op_yVal1(uYc_filtYval1), .op_yVal2(
        uYc_filtYval2), .op_EX_EN(wire_execEnable), .op_DataEN(wire_yAD_Enable), .op_yAddrDiag(uYc_writeDiagAddr), .op_yAddrNonDiag(uYc_writeNonDiagAddr), 
        .op_oneHotDiag(uYc_writeDiagOneHot), .op_oneHotNonDiag(
        uYc_writeNonDiagOneHot) );
  yAddrDecodr unit_yAD1 ( .clock(clock), .reset(reset), .yAD_enable(
        wire_yAD_Enable), .yAD_readRowNum(uYc_opRowNum_from_filtY), 
        .yAD_readRowData(uYc_ySRAM_rowRead1), .yAD_outAddr1(uYc_yMatAddrOut1), 
        .yAD_outAddr2(uYc_yMatAddrOut2), .yAD_dataOutNextCycle(
        wire_dataOuNxtCycle) );
endmodule


module roundRobin ( reset, clock, in_updateYCtrlPathDoneFlag, 
        in_updateYwriteDoneFlag, op_updateYmoduleEnable, op_writeYvalEnable );
  input reset, clock, in_updateYCtrlPathDoneFlag, in_updateYwriteDoneFlag;
  output op_updateYmoduleEnable, op_writeYvalEnable;
  wire   n1, n2, n3, n4, n5, n6;

  DFF_X1 op_updateYmoduleEnable_reg ( .D(n6), .CK(clock), .Q(
        op_updateYmoduleEnable) );
  DFF_X1 op_writeYvalEnable_reg ( .D(n1), .CK(clock), .Q(op_writeYvalEnable)
         );
  NAND2_X2 U4 ( .A1(reset), .A2(n5), .ZN(n6) );
  NAND3_X2 U5 ( .A1(n2), .A2(n3), .A3(op_updateYmoduleEnable), .ZN(n5) );
  INV_X4 U6 ( .A(n4), .ZN(n1) );
  INV_X4 U7 ( .A(in_updateYCtrlPathDoneFlag), .ZN(n2) );
  INV_X4 U8 ( .A(in_updateYwriteDoneFlag), .ZN(n3) );
  OAI211_X2 U3 ( .C1(op_writeYvalEnable), .C2(in_updateYCtrlPathDoneFlag), .A(
        n3), .B(reset), .ZN(n4) );
endmodule


module busArbit ( reset, in_yComputeModuleEnable, in_yWriteModuleEnable, 
        in_controlPathReadAddr1, in_controlPathReadAddr2, in_controlPathWE, 
        in_controlPathWriteAddr, in_controlPathWriteData, 
        in_writePathReadAddr1, in_writePathReadAddr2, in_writePathWE, 
        in_writePathWriteAddr, in_writePathWriteData, op_yReadAddress1, 
        op_yReadAddress2, op_yWriteEnable, op_yWriteAddress, op_writeData );
  input [10:0] in_controlPathReadAddr1;
  input [10:0] in_controlPathReadAddr2;
  input [10:0] in_controlPathWriteAddr;
  input [255:0] in_controlPathWriteData;
  input [10:0] in_writePathReadAddr1;
  input [10:0] in_writePathReadAddr2;
  input [10:0] in_writePathWriteAddr;
  input [255:0] in_writePathWriteData;
  output [10:0] op_yReadAddress1;
  output [10:0] op_yReadAddress2;
  output [10:0] op_yWriteAddress;
  output [255:0] op_writeData;
  input reset, in_yComputeModuleEnable, in_yWriteModuleEnable,
         in_controlPathWE, in_writePathWE;
  output op_yWriteEnable;
  wire   n284, n285, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199;

  INV_X4 U3 ( .A(n285), .ZN(op_yReadAddress1[9]) );
  AOI221_X2 U4 ( .B1(in_controlPathReadAddr1[9]), .B2(n1184), .C1(
        in_writePathReadAddr1[9]), .C2(n1185), .A(n288), .ZN(n285) );
  INV_X4 U5 ( .A(n289), .ZN(op_yReadAddress1[8]) );
  AOI221_X2 U6 ( .B1(in_controlPathReadAddr1[8]), .B2(n1184), .C1(
        in_writePathReadAddr1[8]), .C2(n1185), .A(n288), .ZN(n289) );
  INV_X4 U7 ( .A(n290), .ZN(op_yReadAddress1[7]) );
  AOI221_X2 U8 ( .B1(in_controlPathReadAddr1[7]), .B2(n1184), .C1(
        in_writePathReadAddr1[7]), .C2(n1185), .A(n288), .ZN(n290) );
  INV_X4 U9 ( .A(n291), .ZN(op_yReadAddress1[6]) );
  AOI221_X2 U10 ( .B1(in_controlPathReadAddr1[6]), .B2(n1184), .C1(
        in_writePathReadAddr1[6]), .C2(n1185), .A(n288), .ZN(n291) );
  INV_X4 U11 ( .A(n292), .ZN(op_yReadAddress1[5]) );
  AOI221_X2 U12 ( .B1(in_controlPathReadAddr1[5]), .B2(n1184), .C1(
        in_writePathReadAddr1[5]), .C2(n1185), .A(n288), .ZN(n292) );
  INV_X4 U13 ( .A(n293), .ZN(op_yReadAddress1[4]) );
  AOI221_X2 U14 ( .B1(in_controlPathReadAddr1[4]), .B2(n1184), .C1(
        in_writePathReadAddr1[4]), .C2(n1185), .A(n288), .ZN(n293) );
  INV_X4 U15 ( .A(n294), .ZN(op_yReadAddress1[3]) );
  AOI221_X2 U16 ( .B1(in_controlPathReadAddr1[3]), .B2(n1184), .C1(
        in_writePathReadAddr1[3]), .C2(n1185), .A(n288), .ZN(n294) );
  INV_X4 U17 ( .A(n295), .ZN(op_yReadAddress1[2]) );
  AOI221_X2 U18 ( .B1(in_controlPathReadAddr1[2]), .B2(n1184), .C1(
        in_writePathReadAddr1[2]), .C2(n1185), .A(n288), .ZN(n295) );
  INV_X4 U19 ( .A(n296), .ZN(op_yReadAddress1[10]) );
  AOI221_X2 U20 ( .B1(in_controlPathReadAddr1[10]), .B2(n1184), .C1(
        in_writePathReadAddr1[10]), .C2(n1185), .A(n288), .ZN(n296) );
  INV_X4 U21 ( .A(n297), .ZN(op_yReadAddress1[1]) );
  AOI221_X2 U22 ( .B1(in_controlPathReadAddr1[1]), .B2(n1184), .C1(
        in_writePathReadAddr1[1]), .C2(n1185), .A(n288), .ZN(n297) );
  INV_X4 U23 ( .A(n298), .ZN(op_yReadAddress1[0]) );
  AOI221_X2 U24 ( .B1(in_controlPathReadAddr1[0]), .B2(n1184), .C1(
        in_writePathReadAddr1[0]), .C2(n1185), .A(n1196), .ZN(n298) );
  NAND2_X2 U25 ( .A1(n299), .A2(n300), .ZN(op_yReadAddress2[9]) );
  NAND2_X2 U27 ( .A1(n301), .A2(n300), .ZN(op_yReadAddress2[8]) );
  NAND2_X2 U29 ( .A1(n302), .A2(n300), .ZN(op_yReadAddress2[7]) );
  INV_X4 U31 ( .A(n303), .ZN(op_yReadAddress2[6]) );
  AOI221_X2 U32 ( .B1(in_controlPathReadAddr2[6]), .B2(n1184), .C1(
        in_writePathReadAddr2[6]), .C2(n1185), .A(n1196), .ZN(n303) );
  NAND2_X2 U33 ( .A1(n304), .A2(n300), .ZN(op_yReadAddress2[5]) );
  INV_X4 U35 ( .A(n305), .ZN(op_yReadAddress2[4]) );
  AOI221_X2 U36 ( .B1(in_controlPathReadAddr2[4]), .B2(n1184), .C1(
        in_writePathReadAddr2[4]), .C2(n1185), .A(n1196), .ZN(n305) );
  NAND2_X2 U37 ( .A1(n306), .A2(n300), .ZN(op_yReadAddress2[3]) );
  INV_X4 U39 ( .A(n307), .ZN(op_yReadAddress2[2]) );
  AOI221_X2 U40 ( .B1(in_controlPathReadAddr2[2]), .B2(n1184), .C1(
        in_writePathReadAddr2[2]), .C2(n1185), .A(n1196), .ZN(n307) );
  NAND2_X2 U41 ( .A1(n308), .A2(n300), .ZN(op_yReadAddress2[10]) );
  INV_X4 U43 ( .A(n309), .ZN(op_yReadAddress2[1]) );
  AOI221_X2 U44 ( .B1(in_controlPathReadAddr2[1]), .B2(n1184), .C1(
        in_writePathReadAddr2[1]), .C2(n1185), .A(n1196), .ZN(n309) );
  NAND2_X2 U45 ( .A1(n310), .A2(n300), .ZN(op_yReadAddress2[0]) );
  INV_X4 U47 ( .A(n312), .ZN(op_yWriteEnable) );
  INV_X4 U49 ( .A(n315), .ZN(op_yWriteAddress[9]) );
  AOI221_X2 U50 ( .B1(in_controlPathWriteAddr[9]), .B2(n1184), .C1(
        in_writePathWriteAddr[9]), .C2(n1185), .A(n1196), .ZN(n315) );
  INV_X4 U51 ( .A(n316), .ZN(op_yWriteAddress[8]) );
  AOI221_X2 U52 ( .B1(in_controlPathWriteAddr[8]), .B2(n1184), .C1(
        in_writePathWriteAddr[8]), .C2(n1185), .A(n1196), .ZN(n316) );
  INV_X4 U53 ( .A(n317), .ZN(op_yWriteAddress[7]) );
  AOI221_X2 U54 ( .B1(in_controlPathWriteAddr[7]), .B2(n1184), .C1(
        in_writePathWriteAddr[7]), .C2(n1185), .A(n1196), .ZN(n317) );
  INV_X4 U55 ( .A(n318), .ZN(op_yWriteAddress[6]) );
  AOI221_X2 U56 ( .B1(in_controlPathWriteAddr[6]), .B2(n1184), .C1(
        in_writePathWriteAddr[6]), .C2(n1185), .A(n1196), .ZN(n318) );
  INV_X4 U57 ( .A(n319), .ZN(op_yWriteAddress[5]) );
  AOI221_X2 U58 ( .B1(in_controlPathWriteAddr[5]), .B2(n1184), .C1(
        in_writePathWriteAddr[5]), .C2(n1185), .A(n1196), .ZN(n319) );
  INV_X4 U59 ( .A(n320), .ZN(op_yWriteAddress[4]) );
  AOI221_X2 U60 ( .B1(in_controlPathWriteAddr[4]), .B2(n1184), .C1(
        in_writePathWriteAddr[4]), .C2(n1185), .A(n1196), .ZN(n320) );
  INV_X4 U61 ( .A(n321), .ZN(op_yWriteAddress[3]) );
  AOI221_X2 U62 ( .B1(in_controlPathWriteAddr[3]), .B2(n1184), .C1(
        in_writePathWriteAddr[3]), .C2(n1185), .A(n1196), .ZN(n321) );
  INV_X4 U63 ( .A(n322), .ZN(op_yWriteAddress[2]) );
  AOI221_X2 U64 ( .B1(in_controlPathWriteAddr[2]), .B2(n1184), .C1(
        in_writePathWriteAddr[2]), .C2(n1185), .A(n1196), .ZN(n322) );
  INV_X4 U65 ( .A(n323), .ZN(op_yWriteAddress[10]) );
  AOI221_X2 U66 ( .B1(in_controlPathWriteAddr[10]), .B2(n1184), .C1(
        in_writePathWriteAddr[10]), .C2(n1185), .A(n1196), .ZN(n323) );
  INV_X4 U67 ( .A(n324), .ZN(op_yWriteAddress[1]) );
  AOI221_X2 U68 ( .B1(in_controlPathWriteAddr[1]), .B2(n1184), .C1(
        in_writePathWriteAddr[1]), .C2(n1185), .A(n1196), .ZN(n324) );
  INV_X4 U69 ( .A(n325), .ZN(op_yWriteAddress[0]) );
  AOI221_X2 U70 ( .B1(in_controlPathWriteAddr[0]), .B2(n1184), .C1(
        in_writePathWriteAddr[0]), .C2(n1185), .A(n1196), .ZN(n325) );
  NAND2_X2 U72 ( .A1(in_yWriteModuleEnable), .A2(in_yComputeModuleEnable), 
        .ZN(n311) );
  INV_X4 U73 ( .A(n326), .ZN(op_writeData[99]) );
  INV_X4 U75 ( .A(n327), .ZN(op_writeData[98]) );
  INV_X4 U77 ( .A(n328), .ZN(op_writeData[97]) );
  INV_X4 U79 ( .A(n329), .ZN(op_writeData[96]) );
  INV_X4 U81 ( .A(n330), .ZN(op_writeData[95]) );
  INV_X4 U83 ( .A(n331), .ZN(op_writeData[94]) );
  INV_X4 U85 ( .A(n332), .ZN(op_writeData[93]) );
  INV_X4 U87 ( .A(n333), .ZN(op_writeData[92]) );
  INV_X4 U89 ( .A(n334), .ZN(op_writeData[91]) );
  INV_X4 U91 ( .A(n335), .ZN(op_writeData[90]) );
  INV_X4 U93 ( .A(n336), .ZN(op_writeData[9]) );
  INV_X4 U95 ( .A(n337), .ZN(op_writeData[89]) );
  INV_X4 U97 ( .A(n338), .ZN(op_writeData[88]) );
  INV_X4 U99 ( .A(n339), .ZN(op_writeData[87]) );
  INV_X4 U101 ( .A(n340), .ZN(op_writeData[86]) );
  INV_X4 U103 ( .A(n341), .ZN(op_writeData[85]) );
  INV_X4 U105 ( .A(n342), .ZN(op_writeData[84]) );
  INV_X4 U107 ( .A(n343), .ZN(op_writeData[83]) );
  INV_X4 U109 ( .A(n344), .ZN(op_writeData[82]) );
  INV_X4 U111 ( .A(n345), .ZN(op_writeData[81]) );
  INV_X4 U113 ( .A(n346), .ZN(op_writeData[80]) );
  INV_X4 U115 ( .A(n347), .ZN(op_writeData[8]) );
  INV_X4 U117 ( .A(n348), .ZN(op_writeData[79]) );
  INV_X4 U119 ( .A(n349), .ZN(op_writeData[78]) );
  INV_X4 U121 ( .A(n350), .ZN(op_writeData[77]) );
  INV_X4 U123 ( .A(n351), .ZN(op_writeData[76]) );
  INV_X4 U125 ( .A(n352), .ZN(op_writeData[75]) );
  INV_X4 U127 ( .A(n353), .ZN(op_writeData[74]) );
  INV_X4 U129 ( .A(n354), .ZN(op_writeData[73]) );
  INV_X4 U131 ( .A(n355), .ZN(op_writeData[72]) );
  INV_X4 U133 ( .A(n356), .ZN(op_writeData[71]) );
  INV_X4 U135 ( .A(n357), .ZN(op_writeData[70]) );
  INV_X4 U137 ( .A(n358), .ZN(op_writeData[7]) );
  INV_X4 U139 ( .A(n359), .ZN(op_writeData[69]) );
  INV_X4 U141 ( .A(n360), .ZN(op_writeData[68]) );
  INV_X4 U143 ( .A(n361), .ZN(op_writeData[67]) );
  INV_X4 U145 ( .A(n362), .ZN(op_writeData[66]) );
  INV_X4 U147 ( .A(n363), .ZN(op_writeData[65]) );
  INV_X4 U149 ( .A(n364), .ZN(op_writeData[64]) );
  INV_X4 U151 ( .A(n365), .ZN(op_writeData[63]) );
  INV_X4 U153 ( .A(n366), .ZN(op_writeData[62]) );
  INV_X4 U155 ( .A(n367), .ZN(op_writeData[61]) );
  INV_X4 U157 ( .A(n368), .ZN(op_writeData[60]) );
  INV_X4 U159 ( .A(n369), .ZN(op_writeData[6]) );
  INV_X4 U161 ( .A(n370), .ZN(op_writeData[59]) );
  INV_X4 U163 ( .A(n371), .ZN(op_writeData[58]) );
  INV_X4 U165 ( .A(n372), .ZN(op_writeData[57]) );
  INV_X4 U167 ( .A(n373), .ZN(op_writeData[56]) );
  INV_X4 U169 ( .A(n374), .ZN(op_writeData[55]) );
  INV_X4 U171 ( .A(n375), .ZN(op_writeData[54]) );
  INV_X4 U173 ( .A(n376), .ZN(op_writeData[53]) );
  INV_X4 U175 ( .A(n377), .ZN(op_writeData[52]) );
  INV_X4 U177 ( .A(n378), .ZN(op_writeData[51]) );
  INV_X4 U179 ( .A(n379), .ZN(op_writeData[50]) );
  INV_X4 U181 ( .A(n380), .ZN(op_writeData[5]) );
  INV_X4 U183 ( .A(n381), .ZN(op_writeData[49]) );
  INV_X4 U185 ( .A(n382), .ZN(op_writeData[48]) );
  INV_X4 U187 ( .A(n383), .ZN(op_writeData[47]) );
  INV_X4 U189 ( .A(n384), .ZN(op_writeData[46]) );
  INV_X4 U191 ( .A(n385), .ZN(op_writeData[45]) );
  INV_X4 U193 ( .A(n386), .ZN(op_writeData[44]) );
  INV_X4 U195 ( .A(n387), .ZN(op_writeData[43]) );
  INV_X4 U197 ( .A(n388), .ZN(op_writeData[42]) );
  INV_X4 U199 ( .A(n389), .ZN(op_writeData[41]) );
  INV_X4 U201 ( .A(n390), .ZN(op_writeData[40]) );
  INV_X4 U203 ( .A(n391), .ZN(op_writeData[4]) );
  INV_X4 U205 ( .A(n392), .ZN(op_writeData[39]) );
  INV_X4 U207 ( .A(n393), .ZN(op_writeData[38]) );
  INV_X4 U209 ( .A(n394), .ZN(op_writeData[37]) );
  INV_X4 U211 ( .A(n395), .ZN(op_writeData[36]) );
  INV_X4 U213 ( .A(n396), .ZN(op_writeData[35]) );
  INV_X4 U215 ( .A(n397), .ZN(op_writeData[34]) );
  INV_X4 U217 ( .A(n398), .ZN(op_writeData[33]) );
  INV_X4 U219 ( .A(n399), .ZN(op_writeData[32]) );
  INV_X4 U221 ( .A(n400), .ZN(op_writeData[31]) );
  INV_X4 U223 ( .A(n401), .ZN(op_writeData[30]) );
  INV_X4 U225 ( .A(n402), .ZN(op_writeData[3]) );
  INV_X4 U227 ( .A(n403), .ZN(op_writeData[29]) );
  INV_X4 U229 ( .A(n404), .ZN(op_writeData[28]) );
  INV_X4 U231 ( .A(n405), .ZN(op_writeData[27]) );
  INV_X4 U233 ( .A(n406), .ZN(op_writeData[26]) );
  INV_X4 U235 ( .A(n407), .ZN(op_writeData[255]) );
  INV_X4 U237 ( .A(n408), .ZN(op_writeData[254]) );
  INV_X4 U239 ( .A(n409), .ZN(op_writeData[253]) );
  INV_X4 U241 ( .A(n410), .ZN(op_writeData[252]) );
  INV_X4 U243 ( .A(n411), .ZN(op_writeData[251]) );
  INV_X4 U245 ( .A(n412), .ZN(op_writeData[250]) );
  INV_X4 U247 ( .A(n413), .ZN(op_writeData[25]) );
  INV_X4 U249 ( .A(n414), .ZN(op_writeData[249]) );
  INV_X4 U251 ( .A(n415), .ZN(op_writeData[248]) );
  INV_X4 U253 ( .A(n416), .ZN(op_writeData[247]) );
  INV_X4 U255 ( .A(n417), .ZN(op_writeData[246]) );
  INV_X4 U257 ( .A(n418), .ZN(op_writeData[245]) );
  INV_X4 U259 ( .A(n419), .ZN(op_writeData[244]) );
  INV_X4 U261 ( .A(n420), .ZN(op_writeData[243]) );
  INV_X4 U263 ( .A(n421), .ZN(op_writeData[242]) );
  INV_X4 U265 ( .A(n422), .ZN(op_writeData[241]) );
  INV_X4 U267 ( .A(n423), .ZN(op_writeData[240]) );
  INV_X4 U269 ( .A(n424), .ZN(op_writeData[24]) );
  INV_X4 U271 ( .A(n425), .ZN(op_writeData[239]) );
  INV_X4 U273 ( .A(n426), .ZN(op_writeData[238]) );
  INV_X4 U275 ( .A(n427), .ZN(op_writeData[237]) );
  INV_X4 U277 ( .A(n428), .ZN(op_writeData[236]) );
  INV_X4 U279 ( .A(n429), .ZN(op_writeData[235]) );
  INV_X4 U281 ( .A(n430), .ZN(op_writeData[234]) );
  INV_X4 U283 ( .A(n431), .ZN(op_writeData[233]) );
  INV_X4 U285 ( .A(n432), .ZN(op_writeData[232]) );
  INV_X4 U287 ( .A(n433), .ZN(op_writeData[231]) );
  INV_X4 U289 ( .A(n434), .ZN(op_writeData[230]) );
  INV_X4 U291 ( .A(n435), .ZN(op_writeData[23]) );
  INV_X4 U293 ( .A(n436), .ZN(op_writeData[229]) );
  INV_X4 U295 ( .A(n437), .ZN(op_writeData[228]) );
  INV_X4 U297 ( .A(n438), .ZN(op_writeData[227]) );
  INV_X4 U299 ( .A(n439), .ZN(op_writeData[226]) );
  INV_X4 U301 ( .A(n440), .ZN(op_writeData[225]) );
  INV_X4 U303 ( .A(n441), .ZN(op_writeData[224]) );
  INV_X4 U305 ( .A(n442), .ZN(op_writeData[223]) );
  INV_X4 U307 ( .A(n443), .ZN(op_writeData[222]) );
  INV_X4 U309 ( .A(n444), .ZN(op_writeData[221]) );
  INV_X4 U311 ( .A(n445), .ZN(op_writeData[220]) );
  INV_X4 U313 ( .A(n446), .ZN(op_writeData[22]) );
  INV_X4 U315 ( .A(n447), .ZN(op_writeData[219]) );
  INV_X4 U317 ( .A(n448), .ZN(op_writeData[218]) );
  INV_X4 U319 ( .A(n449), .ZN(op_writeData[217]) );
  INV_X4 U321 ( .A(n450), .ZN(op_writeData[216]) );
  INV_X4 U323 ( .A(n451), .ZN(op_writeData[215]) );
  INV_X4 U325 ( .A(n452), .ZN(op_writeData[214]) );
  INV_X4 U327 ( .A(n453), .ZN(op_writeData[213]) );
  INV_X4 U329 ( .A(n454), .ZN(op_writeData[212]) );
  INV_X4 U331 ( .A(n455), .ZN(op_writeData[211]) );
  INV_X4 U333 ( .A(n456), .ZN(op_writeData[210]) );
  INV_X4 U335 ( .A(n457), .ZN(op_writeData[21]) );
  INV_X4 U337 ( .A(n458), .ZN(op_writeData[209]) );
  INV_X4 U339 ( .A(n459), .ZN(op_writeData[208]) );
  INV_X4 U341 ( .A(n460), .ZN(op_writeData[207]) );
  INV_X4 U343 ( .A(n461), .ZN(op_writeData[206]) );
  INV_X4 U345 ( .A(n462), .ZN(op_writeData[205]) );
  INV_X4 U347 ( .A(n463), .ZN(op_writeData[204]) );
  INV_X4 U349 ( .A(n464), .ZN(op_writeData[203]) );
  INV_X4 U351 ( .A(n465), .ZN(op_writeData[202]) );
  INV_X4 U353 ( .A(n466), .ZN(op_writeData[201]) );
  INV_X4 U355 ( .A(n467), .ZN(op_writeData[200]) );
  INV_X4 U357 ( .A(n468), .ZN(op_writeData[20]) );
  INV_X4 U359 ( .A(n469), .ZN(op_writeData[2]) );
  INV_X4 U361 ( .A(n470), .ZN(op_writeData[199]) );
  INV_X4 U363 ( .A(n471), .ZN(op_writeData[198]) );
  INV_X4 U365 ( .A(n472), .ZN(op_writeData[197]) );
  INV_X4 U367 ( .A(n473), .ZN(op_writeData[196]) );
  INV_X4 U369 ( .A(n474), .ZN(op_writeData[195]) );
  INV_X4 U371 ( .A(n475), .ZN(op_writeData[194]) );
  INV_X4 U373 ( .A(n476), .ZN(op_writeData[193]) );
  INV_X4 U375 ( .A(n477), .ZN(op_writeData[192]) );
  INV_X4 U377 ( .A(n478), .ZN(op_writeData[191]) );
  INV_X4 U379 ( .A(n479), .ZN(op_writeData[190]) );
  INV_X4 U381 ( .A(n480), .ZN(op_writeData[19]) );
  INV_X4 U383 ( .A(n481), .ZN(op_writeData[189]) );
  INV_X4 U385 ( .A(n482), .ZN(op_writeData[188]) );
  INV_X4 U387 ( .A(n483), .ZN(op_writeData[187]) );
  INV_X4 U389 ( .A(n484), .ZN(op_writeData[186]) );
  INV_X4 U391 ( .A(n485), .ZN(op_writeData[185]) );
  INV_X4 U393 ( .A(n486), .ZN(op_writeData[184]) );
  INV_X4 U395 ( .A(n487), .ZN(op_writeData[183]) );
  INV_X4 U397 ( .A(n488), .ZN(op_writeData[182]) );
  INV_X4 U399 ( .A(n489), .ZN(op_writeData[181]) );
  INV_X4 U401 ( .A(n490), .ZN(op_writeData[180]) );
  INV_X4 U403 ( .A(n491), .ZN(op_writeData[18]) );
  INV_X4 U405 ( .A(n492), .ZN(op_writeData[179]) );
  INV_X4 U407 ( .A(n493), .ZN(op_writeData[178]) );
  INV_X4 U409 ( .A(n494), .ZN(op_writeData[177]) );
  INV_X4 U411 ( .A(n495), .ZN(op_writeData[176]) );
  INV_X4 U413 ( .A(n496), .ZN(op_writeData[175]) );
  INV_X4 U415 ( .A(n497), .ZN(op_writeData[174]) );
  INV_X4 U417 ( .A(n498), .ZN(op_writeData[173]) );
  INV_X4 U419 ( .A(n499), .ZN(op_writeData[172]) );
  INV_X4 U421 ( .A(n500), .ZN(op_writeData[171]) );
  INV_X4 U423 ( .A(n501), .ZN(op_writeData[170]) );
  INV_X4 U425 ( .A(n502), .ZN(op_writeData[17]) );
  INV_X4 U427 ( .A(n503), .ZN(op_writeData[169]) );
  INV_X4 U429 ( .A(n504), .ZN(op_writeData[168]) );
  INV_X4 U431 ( .A(n505), .ZN(op_writeData[167]) );
  INV_X4 U433 ( .A(n506), .ZN(op_writeData[166]) );
  INV_X4 U435 ( .A(n507), .ZN(op_writeData[165]) );
  INV_X4 U437 ( .A(n508), .ZN(op_writeData[164]) );
  INV_X4 U439 ( .A(n509), .ZN(op_writeData[163]) );
  INV_X4 U441 ( .A(n510), .ZN(op_writeData[162]) );
  INV_X4 U443 ( .A(n511), .ZN(op_writeData[161]) );
  INV_X4 U445 ( .A(n512), .ZN(op_writeData[160]) );
  INV_X4 U447 ( .A(n513), .ZN(op_writeData[16]) );
  INV_X4 U449 ( .A(n514), .ZN(op_writeData[159]) );
  INV_X4 U451 ( .A(n515), .ZN(op_writeData[158]) );
  INV_X4 U453 ( .A(n516), .ZN(op_writeData[157]) );
  INV_X4 U455 ( .A(n517), .ZN(op_writeData[156]) );
  INV_X4 U457 ( .A(n518), .ZN(op_writeData[155]) );
  INV_X4 U459 ( .A(n519), .ZN(op_writeData[154]) );
  INV_X4 U461 ( .A(n520), .ZN(op_writeData[153]) );
  INV_X4 U463 ( .A(n521), .ZN(op_writeData[152]) );
  INV_X4 U465 ( .A(n522), .ZN(op_writeData[151]) );
  INV_X4 U467 ( .A(n523), .ZN(op_writeData[150]) );
  INV_X4 U469 ( .A(n524), .ZN(op_writeData[15]) );
  INV_X4 U471 ( .A(n525), .ZN(op_writeData[149]) );
  INV_X4 U473 ( .A(n526), .ZN(op_writeData[148]) );
  INV_X4 U475 ( .A(n527), .ZN(op_writeData[147]) );
  INV_X4 U477 ( .A(n528), .ZN(op_writeData[146]) );
  INV_X4 U479 ( .A(n529), .ZN(op_writeData[145]) );
  INV_X4 U481 ( .A(n530), .ZN(op_writeData[144]) );
  INV_X4 U483 ( .A(n531), .ZN(op_writeData[143]) );
  INV_X4 U485 ( .A(n532), .ZN(op_writeData[142]) );
  INV_X4 U487 ( .A(n533), .ZN(op_writeData[141]) );
  INV_X4 U489 ( .A(n534), .ZN(op_writeData[140]) );
  INV_X4 U491 ( .A(n535), .ZN(op_writeData[14]) );
  INV_X4 U493 ( .A(n536), .ZN(op_writeData[139]) );
  INV_X4 U495 ( .A(n537), .ZN(op_writeData[138]) );
  INV_X4 U497 ( .A(n538), .ZN(op_writeData[137]) );
  INV_X4 U499 ( .A(n539), .ZN(op_writeData[136]) );
  INV_X4 U501 ( .A(n540), .ZN(op_writeData[135]) );
  INV_X4 U503 ( .A(n541), .ZN(op_writeData[134]) );
  INV_X4 U505 ( .A(n542), .ZN(op_writeData[133]) );
  INV_X4 U507 ( .A(n543), .ZN(op_writeData[132]) );
  INV_X4 U509 ( .A(n544), .ZN(op_writeData[131]) );
  INV_X4 U511 ( .A(n545), .ZN(op_writeData[130]) );
  INV_X4 U513 ( .A(n546), .ZN(op_writeData[13]) );
  INV_X4 U515 ( .A(n547), .ZN(op_writeData[129]) );
  INV_X4 U517 ( .A(n548), .ZN(op_writeData[128]) );
  INV_X4 U519 ( .A(n549), .ZN(op_writeData[127]) );
  INV_X4 U521 ( .A(n550), .ZN(op_writeData[126]) );
  INV_X4 U523 ( .A(n551), .ZN(op_writeData[125]) );
  INV_X4 U525 ( .A(n552), .ZN(op_writeData[124]) );
  INV_X4 U527 ( .A(n553), .ZN(op_writeData[123]) );
  INV_X4 U529 ( .A(n554), .ZN(op_writeData[122]) );
  INV_X4 U531 ( .A(n555), .ZN(op_writeData[121]) );
  INV_X4 U533 ( .A(n556), .ZN(op_writeData[120]) );
  INV_X4 U535 ( .A(n557), .ZN(op_writeData[12]) );
  INV_X4 U537 ( .A(n558), .ZN(op_writeData[119]) );
  INV_X4 U539 ( .A(n559), .ZN(op_writeData[118]) );
  INV_X4 U541 ( .A(n560), .ZN(op_writeData[117]) );
  INV_X4 U543 ( .A(n561), .ZN(op_writeData[116]) );
  INV_X4 U545 ( .A(n562), .ZN(op_writeData[115]) );
  INV_X4 U547 ( .A(n563), .ZN(op_writeData[114]) );
  INV_X4 U549 ( .A(n564), .ZN(op_writeData[113]) );
  INV_X4 U551 ( .A(n565), .ZN(op_writeData[112]) );
  INV_X4 U553 ( .A(n566), .ZN(op_writeData[111]) );
  INV_X4 U555 ( .A(n567), .ZN(op_writeData[110]) );
  INV_X4 U557 ( .A(n568), .ZN(op_writeData[11]) );
  INV_X4 U559 ( .A(n569), .ZN(op_writeData[109]) );
  INV_X4 U561 ( .A(n570), .ZN(op_writeData[108]) );
  INV_X4 U563 ( .A(n571), .ZN(op_writeData[107]) );
  INV_X4 U565 ( .A(n572), .ZN(op_writeData[106]) );
  INV_X4 U567 ( .A(n573), .ZN(op_writeData[105]) );
  INV_X4 U569 ( .A(n574), .ZN(op_writeData[104]) );
  INV_X4 U571 ( .A(n575), .ZN(op_writeData[103]) );
  INV_X4 U573 ( .A(n576), .ZN(op_writeData[102]) );
  INV_X4 U575 ( .A(n577), .ZN(op_writeData[101]) );
  INV_X4 U577 ( .A(n578), .ZN(op_writeData[100]) );
  INV_X4 U579 ( .A(n579), .ZN(op_writeData[10]) );
  INV_X4 U581 ( .A(n580), .ZN(op_writeData[1]) );
  INV_X4 U583 ( .A(n581), .ZN(op_writeData[0]) );
  INV_X4 U586 ( .A(in_yComputeModuleEnable), .ZN(n284) );
  AND2_X1 U587 ( .A1(reset), .A2(n311), .ZN(n300) );
  AND2_X4 U26 ( .A1(n1184), .A2(reset), .ZN(n313) );
  AND2_X4 U28 ( .A1(n1185), .A2(reset), .ZN(n1183) );
  NOR2_X4 U30 ( .A1(n284), .A2(in_yWriteModuleEnable), .ZN(n1184) );
  AND2_X4 U34 ( .A1(in_yWriteModuleEnable), .A2(n284), .ZN(n1185) );
  INV_X4 U80 ( .A(n1199), .ZN(n1190) );
  INV_X4 U82 ( .A(n313), .ZN(n1195) );
  INV_X4 U84 ( .A(n1197), .ZN(n1196) );
  AOI22_X2 U86 ( .A1(in_controlPathWriteData[0]), .A2(n313), .B1(
        in_writePathWriteData[0]), .B2(n1186), .ZN(n581) );
  AOI22_X2 U88 ( .A1(in_controlPathWriteData[1]), .A2(n1192), .B1(
        in_writePathWriteData[1]), .B2(n1187), .ZN(n580) );
  AOI22_X2 U90 ( .A1(in_controlPathWriteData[2]), .A2(n1192), .B1(
        in_writePathWriteData[2]), .B2(n1189), .ZN(n469) );
  AOI22_X2 U92 ( .A1(in_controlPathWriteData[3]), .A2(n313), .B1(
        in_writePathWriteData[3]), .B2(n1187), .ZN(n402) );
  AOI22_X2 U94 ( .A1(in_controlPathWriteData[4]), .A2(n313), .B1(
        in_writePathWriteData[4]), .B2(n1188), .ZN(n391) );
  AOI22_X2 U96 ( .A1(in_controlPathWriteData[5]), .A2(n1194), .B1(
        in_writePathWriteData[5]), .B2(n1189), .ZN(n380) );
  AOI22_X2 U98 ( .A1(in_controlPathWriteData[6]), .A2(n1193), .B1(
        in_writePathWriteData[6]), .B2(n1186), .ZN(n369) );
  AOI22_X2 U100 ( .A1(in_controlPathWriteData[7]), .A2(n313), .B1(
        in_writePathWriteData[7]), .B2(n1188), .ZN(n358) );
  AOI22_X2 U102 ( .A1(in_controlPathWriteData[8]), .A2(n1194), .B1(
        in_writePathWriteData[8]), .B2(n1187), .ZN(n347) );
  AOI22_X2 U104 ( .A1(in_controlPathWriteData[9]), .A2(n1191), .B1(
        in_writePathWriteData[9]), .B2(n1186), .ZN(n336) );
  AOI22_X2 U106 ( .A1(in_controlPathWriteData[10]), .A2(n1193), .B1(
        in_writePathWriteData[10]), .B2(n1186), .ZN(n579) );
  AOI22_X2 U108 ( .A1(in_controlPathWriteData[11]), .A2(n1194), .B1(
        in_writePathWriteData[11]), .B2(n1187), .ZN(n568) );
  AOI22_X2 U110 ( .A1(in_controlPathWriteData[12]), .A2(n1191), .B1(
        in_writePathWriteData[12]), .B2(n1199), .ZN(n557) );
  AOI22_X2 U112 ( .A1(in_controlPathWriteData[13]), .A2(n1192), .B1(
        in_writePathWriteData[13]), .B2(n1199), .ZN(n546) );
  AOI22_X2 U114 ( .A1(in_controlPathWriteData[14]), .A2(n313), .B1(
        in_writePathWriteData[14]), .B2(n1189), .ZN(n535) );
  AOI22_X2 U116 ( .A1(in_controlPathWriteData[15]), .A2(n1194), .B1(
        in_writePathWriteData[15]), .B2(n1187), .ZN(n524) );
  AOI22_X2 U118 ( .A1(in_controlPathWriteData[16]), .A2(n1192), .B1(
        in_writePathWriteData[16]), .B2(n1189), .ZN(n513) );
  AOI22_X2 U120 ( .A1(in_controlPathWriteData[17]), .A2(n1193), .B1(
        in_writePathWriteData[17]), .B2(n1199), .ZN(n502) );
  AOI22_X2 U122 ( .A1(in_controlPathWriteData[18]), .A2(n1191), .B1(
        in_writePathWriteData[18]), .B2(n1189), .ZN(n491) );
  AOI22_X2 U124 ( .A1(in_controlPathWriteData[19]), .A2(n1194), .B1(
        in_writePathWriteData[19]), .B2(n1188), .ZN(n480) );
  AOI22_X2 U126 ( .A1(in_controlPathWriteData[20]), .A2(n1193), .B1(
        in_writePathWriteData[20]), .B2(n1188), .ZN(n468) );
  AOI22_X2 U128 ( .A1(in_controlPathWriteData[21]), .A2(n313), .B1(
        in_writePathWriteData[21]), .B2(n1186), .ZN(n457) );
  AOI22_X2 U130 ( .A1(in_controlPathWriteData[22]), .A2(n1191), .B1(
        in_writePathWriteData[22]), .B2(n1189), .ZN(n446) );
  AOI22_X2 U132 ( .A1(in_controlPathWriteData[23]), .A2(n313), .B1(
        in_writePathWriteData[23]), .B2(n1188), .ZN(n435) );
  AOI22_X2 U134 ( .A1(in_controlPathWriteData[24]), .A2(n1192), .B1(
        in_writePathWriteData[24]), .B2(n1186), .ZN(n424) );
  AOI22_X2 U136 ( .A1(in_controlPathWriteData[25]), .A2(n1192), .B1(
        in_writePathWriteData[25]), .B2(n1188), .ZN(n413) );
  AOI22_X2 U138 ( .A1(in_controlPathWriteData[26]), .A2(n1194), .B1(
        in_writePathWriteData[26]), .B2(n1187), .ZN(n406) );
  AOI22_X2 U140 ( .A1(in_controlPathWriteData[27]), .A2(n313), .B1(
        in_writePathWriteData[27]), .B2(n1199), .ZN(n405) );
  AOI22_X2 U142 ( .A1(in_controlPathWriteData[28]), .A2(n1191), .B1(
        in_writePathWriteData[28]), .B2(n1199), .ZN(n404) );
  AOI22_X2 U144 ( .A1(in_controlPathWriteData[29]), .A2(n1193), .B1(
        in_writePathWriteData[29]), .B2(n1199), .ZN(n403) );
  AOI22_X2 U146 ( .A1(in_controlPathWriteData[30]), .A2(n1191), .B1(
        in_writePathWriteData[30]), .B2(n1186), .ZN(n401) );
  AOI22_X2 U148 ( .A1(in_controlPathWriteData[31]), .A2(n1192), .B1(
        in_writePathWriteData[31]), .B2(n1186), .ZN(n400) );
  AOI22_X2 U150 ( .A1(in_controlPathWriteData[32]), .A2(n313), .B1(
        in_writePathWriteData[32]), .B2(n1187), .ZN(n399) );
  AOI22_X2 U152 ( .A1(in_controlPathWriteData[33]), .A2(n313), .B1(
        in_writePathWriteData[33]), .B2(n1189), .ZN(n398) );
  AOI22_X2 U154 ( .A1(in_controlPathWriteData[34]), .A2(n313), .B1(
        in_writePathWriteData[34]), .B2(n1187), .ZN(n397) );
  AOI22_X2 U156 ( .A1(in_controlPathWriteData[35]), .A2(n313), .B1(
        in_writePathWriteData[35]), .B2(n1189), .ZN(n396) );
  AOI22_X2 U158 ( .A1(in_controlPathWriteData[36]), .A2(n1193), .B1(
        in_writePathWriteData[36]), .B2(n1187), .ZN(n395) );
  AOI22_X2 U160 ( .A1(in_controlPathWriteData[37]), .A2(n1192), .B1(
        in_writePathWriteData[37]), .B2(n1189), .ZN(n394) );
  AOI22_X2 U162 ( .A1(in_controlPathWriteData[38]), .A2(n1194), .B1(
        in_writePathWriteData[38]), .B2(n1188), .ZN(n393) );
  AOI22_X2 U164 ( .A1(in_controlPathWriteData[39]), .A2(n1194), .B1(
        in_writePathWriteData[39]), .B2(n1188), .ZN(n392) );
  AOI22_X2 U166 ( .A1(in_controlPathWriteData[40]), .A2(n1193), .B1(
        in_writePathWriteData[40]), .B2(n1188), .ZN(n390) );
  AOI22_X2 U168 ( .A1(in_controlPathWriteData[41]), .A2(n1193), .B1(
        in_writePathWriteData[41]), .B2(n1186), .ZN(n389) );
  AOI22_X2 U170 ( .A1(in_controlPathWriteData[42]), .A2(n1194), .B1(
        in_writePathWriteData[42]), .B2(n1186), .ZN(n388) );
  AOI22_X2 U172 ( .A1(in_controlPathWriteData[43]), .A2(n1191), .B1(
        in_writePathWriteData[43]), .B2(n1187), .ZN(n387) );
  AOI22_X2 U174 ( .A1(in_controlPathWriteData[44]), .A2(n1192), .B1(
        in_writePathWriteData[44]), .B2(n1189), .ZN(n386) );
  AOI22_X2 U176 ( .A1(in_controlPathWriteData[45]), .A2(n1193), .B1(
        in_writePathWriteData[45]), .B2(n1189), .ZN(n385) );
  AOI22_X2 U178 ( .A1(in_controlPathWriteData[46]), .A2(n1194), .B1(
        in_writePathWriteData[46]), .B2(n1186), .ZN(n384) );
  AOI22_X2 U180 ( .A1(in_controlPathWriteData[47]), .A2(n1191), .B1(
        in_writePathWriteData[47]), .B2(n1187), .ZN(n383) );
  AOI22_X2 U182 ( .A1(in_controlPathWriteData[48]), .A2(n1192), .B1(
        in_writePathWriteData[48]), .B2(n1188), .ZN(n382) );
  AOI22_X2 U184 ( .A1(in_controlPathWriteData[49]), .A2(n1193), .B1(
        in_writePathWriteData[49]), .B2(n1187), .ZN(n381) );
  AOI22_X2 U186 ( .A1(in_controlPathWriteData[50]), .A2(n1194), .B1(
        in_writePathWriteData[50]), .B2(n1188), .ZN(n379) );
  AOI22_X2 U188 ( .A1(in_controlPathWriteData[51]), .A2(n1191), .B1(
        in_writePathWriteData[51]), .B2(n1189), .ZN(n378) );
  AOI22_X2 U190 ( .A1(in_controlPathWriteData[52]), .A2(n1191), .B1(
        in_writePathWriteData[52]), .B2(n1186), .ZN(n377) );
  AOI22_X2 U192 ( .A1(in_controlPathWriteData[53]), .A2(n1192), .B1(
        in_writePathWriteData[53]), .B2(n1186), .ZN(n376) );
  AOI22_X2 U194 ( .A1(in_controlPathWriteData[54]), .A2(n1193), .B1(
        in_writePathWriteData[54]), .B2(n1199), .ZN(n375) );
  AOI22_X2 U196 ( .A1(in_controlPathWriteData[55]), .A2(n1194), .B1(
        in_writePathWriteData[55]), .B2(n1199), .ZN(n374) );
  AOI22_X2 U198 ( .A1(in_controlPathWriteData[56]), .A2(n1191), .B1(
        in_writePathWriteData[56]), .B2(n1199), .ZN(n373) );
  AOI22_X2 U200 ( .A1(in_controlPathWriteData[57]), .A2(n1192), .B1(
        in_writePathWriteData[57]), .B2(n1199), .ZN(n372) );
  AOI22_X2 U202 ( .A1(in_controlPathWriteData[58]), .A2(n1193), .B1(
        in_writePathWriteData[58]), .B2(n1199), .ZN(n371) );
  AOI22_X2 U204 ( .A1(in_controlPathWriteData[59]), .A2(n1194), .B1(
        in_writePathWriteData[59]), .B2(n1199), .ZN(n370) );
  AOI22_X2 U206 ( .A1(in_controlPathWriteData[60]), .A2(n1191), .B1(
        in_writePathWriteData[60]), .B2(n1199), .ZN(n368) );
  AOI22_X2 U208 ( .A1(in_controlPathWriteData[61]), .A2(n1192), .B1(
        in_writePathWriteData[61]), .B2(n1199), .ZN(n367) );
  AOI22_X2 U210 ( .A1(in_controlPathWriteData[62]), .A2(n1193), .B1(
        in_writePathWriteData[62]), .B2(n1199), .ZN(n366) );
  AOI22_X2 U212 ( .A1(in_controlPathWriteData[63]), .A2(n313), .B1(
        in_writePathWriteData[63]), .B2(n1188), .ZN(n365) );
  AOI22_X2 U214 ( .A1(in_controlPathWriteData[64]), .A2(n313), .B1(
        in_writePathWriteData[64]), .B2(n1187), .ZN(n364) );
  AOI22_X2 U216 ( .A1(in_controlPathWriteData[65]), .A2(n313), .B1(
        in_writePathWriteData[65]), .B2(n1189), .ZN(n363) );
  AOI22_X2 U218 ( .A1(in_controlPathWriteData[66]), .A2(n313), .B1(
        in_writePathWriteData[66]), .B2(n1187), .ZN(n362) );
  AOI22_X2 U220 ( .A1(in_controlPathWriteData[67]), .A2(n313), .B1(
        in_writePathWriteData[67]), .B2(n1188), .ZN(n361) );
  AOI22_X2 U222 ( .A1(in_controlPathWriteData[68]), .A2(n313), .B1(
        in_writePathWriteData[68]), .B2(n1189), .ZN(n360) );
  AOI22_X2 U224 ( .A1(in_controlPathWriteData[69]), .A2(n313), .B1(
        in_writePathWriteData[69]), .B2(n1186), .ZN(n359) );
  AOI22_X2 U226 ( .A1(in_controlPathWriteData[70]), .A2(n313), .B1(
        in_writePathWriteData[70]), .B2(n1187), .ZN(n357) );
  AOI22_X2 U228 ( .A1(in_controlPathWriteData[71]), .A2(n313), .B1(
        in_writePathWriteData[71]), .B2(n1199), .ZN(n356) );
  AOI22_X2 U230 ( .A1(in_controlPathWriteData[72]), .A2(n313), .B1(
        in_writePathWriteData[72]), .B2(n1199), .ZN(n355) );
  AOI22_X2 U232 ( .A1(in_controlPathWriteData[73]), .A2(n313), .B1(
        in_writePathWriteData[73]), .B2(n1188), .ZN(n354) );
  AOI22_X2 U234 ( .A1(in_controlPathWriteData[74]), .A2(n1194), .B1(
        in_writePathWriteData[74]), .B2(n1186), .ZN(n353) );
  AOI22_X2 U236 ( .A1(in_controlPathWriteData[75]), .A2(n1191), .B1(
        in_writePathWriteData[75]), .B2(n1186), .ZN(n352) );
  AOI22_X2 U238 ( .A1(in_controlPathWriteData[76]), .A2(n1192), .B1(
        in_writePathWriteData[76]), .B2(n1189), .ZN(n351) );
  AOI22_X2 U240 ( .A1(in_controlPathWriteData[77]), .A2(n1193), .B1(
        in_writePathWriteData[77]), .B2(n1188), .ZN(n350) );
  AOI22_X2 U242 ( .A1(in_controlPathWriteData[78]), .A2(n1194), .B1(
        in_writePathWriteData[78]), .B2(n1187), .ZN(n349) );
  AOI22_X2 U244 ( .A1(in_controlPathWriteData[79]), .A2(n1191), .B1(
        in_writePathWriteData[79]), .B2(n1199), .ZN(n348) );
  AOI22_X2 U246 ( .A1(in_controlPathWriteData[80]), .A2(n1192), .B1(
        in_writePathWriteData[80]), .B2(n1199), .ZN(n346) );
  AOI22_X2 U248 ( .A1(in_controlPathWriteData[81]), .A2(n1193), .B1(
        in_writePathWriteData[81]), .B2(n1199), .ZN(n345) );
  AOI22_X2 U250 ( .A1(in_controlPathWriteData[82]), .A2(n1194), .B1(
        in_writePathWriteData[82]), .B2(n1199), .ZN(n344) );
  AOI22_X2 U252 ( .A1(in_controlPathWriteData[83]), .A2(n1191), .B1(
        in_writePathWriteData[83]), .B2(n1199), .ZN(n343) );
  AOI22_X2 U254 ( .A1(in_controlPathWriteData[84]), .A2(n1192), .B1(
        in_writePathWriteData[84]), .B2(n1199), .ZN(n342) );
  AOI22_X2 U256 ( .A1(in_controlPathWriteData[85]), .A2(n1191), .B1(
        in_writePathWriteData[85]), .B2(n1187), .ZN(n341) );
  AOI22_X2 U258 ( .A1(in_controlPathWriteData[86]), .A2(n1192), .B1(
        in_writePathWriteData[86]), .B2(n1189), .ZN(n340) );
  AOI22_X2 U260 ( .A1(in_controlPathWriteData[87]), .A2(n1194), .B1(
        in_writePathWriteData[87]), .B2(n1188), .ZN(n339) );
  AOI22_X2 U262 ( .A1(in_controlPathWriteData[88]), .A2(n313), .B1(
        in_writePathWriteData[88]), .B2(n1186), .ZN(n338) );
  AOI22_X2 U264 ( .A1(in_controlPathWriteData[89]), .A2(n1193), .B1(
        in_writePathWriteData[89]), .B2(n1187), .ZN(n337) );
  AOI22_X2 U266 ( .A1(in_controlPathWriteData[90]), .A2(n1191), .B1(
        in_writePathWriteData[90]), .B2(n1189), .ZN(n335) );
  AOI22_X2 U268 ( .A1(in_controlPathWriteData[91]), .A2(n1192), .B1(
        in_writePathWriteData[91]), .B2(n1188), .ZN(n334) );
  AOI22_X2 U270 ( .A1(in_controlPathWriteData[92]), .A2(n1193), .B1(
        in_writePathWriteData[92]), .B2(n1186), .ZN(n333) );
  AOI22_X2 U272 ( .A1(in_controlPathWriteData[93]), .A2(n313), .B1(
        in_writePathWriteData[93]), .B2(n1187), .ZN(n332) );
  AOI22_X2 U274 ( .A1(in_controlPathWriteData[94]), .A2(n1192), .B1(
        in_writePathWriteData[94]), .B2(n1189), .ZN(n331) );
  AOI22_X2 U276 ( .A1(in_controlPathWriteData[95]), .A2(n1193), .B1(
        in_writePathWriteData[95]), .B2(n1188), .ZN(n330) );
  AOI22_X2 U278 ( .A1(in_controlPathWriteData[100]), .A2(n1194), .B1(
        in_writePathWriteData[100]), .B2(n1186), .ZN(n578) );
  AOI22_X2 U280 ( .A1(in_controlPathWriteData[101]), .A2(n1194), .B1(
        in_writePathWriteData[101]), .B2(n1187), .ZN(n577) );
  AOI22_X2 U282 ( .A1(in_controlPathWriteData[102]), .A2(n1193), .B1(
        in_writePathWriteData[102]), .B2(n1189), .ZN(n576) );
  AOI22_X2 U284 ( .A1(in_controlPathWriteData[103]), .A2(n1191), .B1(
        in_writePathWriteData[103]), .B2(n1186), .ZN(n575) );
  AOI22_X2 U286 ( .A1(in_controlPathWriteData[104]), .A2(n1194), .B1(
        in_writePathWriteData[104]), .B2(n1189), .ZN(n574) );
  AOI22_X2 U288 ( .A1(in_controlPathWriteData[105]), .A2(n1191), .B1(
        in_writePathWriteData[105]), .B2(n1189), .ZN(n573) );
  AOI22_X2 U290 ( .A1(in_controlPathWriteData[106]), .A2(n1191), .B1(
        in_writePathWriteData[106]), .B2(n1188), .ZN(n572) );
  AOI22_X2 U292 ( .A1(in_controlPathWriteData[107]), .A2(n313), .B1(
        in_writePathWriteData[107]), .B2(n1188), .ZN(n571) );
  AOI22_X2 U294 ( .A1(in_controlPathWriteData[108]), .A2(n1194), .B1(
        in_writePathWriteData[108]), .B2(n1186), .ZN(n570) );
  AOI22_X2 U296 ( .A1(in_controlPathWriteData[109]), .A2(n1191), .B1(
        in_writePathWriteData[109]), .B2(n1186), .ZN(n569) );
  AOI22_X2 U298 ( .A1(in_controlPathWriteData[110]), .A2(n1192), .B1(
        in_writePathWriteData[110]), .B2(n1188), .ZN(n567) );
  AOI22_X2 U300 ( .A1(in_controlPathWriteData[111]), .A2(n1193), .B1(
        in_writePathWriteData[111]), .B2(n1186), .ZN(n566) );
  AOI22_X2 U302 ( .A1(in_controlPathWriteData[112]), .A2(n1194), .B1(
        in_writePathWriteData[112]), .B2(n1199), .ZN(n565) );
  AOI22_X2 U304 ( .A1(in_controlPathWriteData[113]), .A2(n1191), .B1(
        in_writePathWriteData[113]), .B2(n1199), .ZN(n564) );
  AOI22_X2 U306 ( .A1(in_controlPathWriteData[114]), .A2(n1192), .B1(
        in_writePathWriteData[114]), .B2(n1187), .ZN(n563) );
  AOI22_X2 U308 ( .A1(in_controlPathWriteData[115]), .A2(n1193), .B1(
        in_writePathWriteData[115]), .B2(n1187), .ZN(n562) );
  AOI22_X2 U310 ( .A1(in_controlPathWriteData[116]), .A2(n1194), .B1(
        in_writePathWriteData[116]), .B2(n1189), .ZN(n561) );
  AOI22_X2 U312 ( .A1(in_controlPathWriteData[117]), .A2(n1191), .B1(
        in_writePathWriteData[117]), .B2(n1189), .ZN(n560) );
  AOI22_X2 U314 ( .A1(in_controlPathWriteData[118]), .A2(n1192), .B1(
        in_writePathWriteData[118]), .B2(n1188), .ZN(n559) );
  AOI22_X2 U316 ( .A1(in_controlPathWriteData[119]), .A2(n1193), .B1(
        in_writePathWriteData[119]), .B2(n1186), .ZN(n558) );
  AOI22_X2 U318 ( .A1(in_controlPathWriteData[120]), .A2(n1192), .B1(
        in_writePathWriteData[120]), .B2(n1187), .ZN(n556) );
  AOI22_X2 U320 ( .A1(in_controlPathWriteData[121]), .A2(n1194), .B1(
        in_writePathWriteData[121]), .B2(n1189), .ZN(n555) );
  AOI22_X2 U322 ( .A1(in_controlPathWriteData[122]), .A2(n1191), .B1(
        in_writePathWriteData[122]), .B2(n1188), .ZN(n554) );
  AOI22_X2 U324 ( .A1(in_controlPathWriteData[123]), .A2(n1193), .B1(
        in_writePathWriteData[123]), .B2(n1199), .ZN(n553) );
  AOI22_X2 U326 ( .A1(in_controlPathWriteData[124]), .A2(n1192), .B1(
        in_writePathWriteData[124]), .B2(n1199), .ZN(n552) );
  AOI22_X2 U328 ( .A1(in_controlPathWriteData[125]), .A2(n1194), .B1(
        in_writePathWriteData[125]), .B2(n1187), .ZN(n551) );
  AOI22_X2 U330 ( .A1(in_controlPathWriteData[126]), .A2(n1191), .B1(
        in_writePathWriteData[126]), .B2(n1189), .ZN(n550) );
  AOI22_X2 U332 ( .A1(in_controlPathWriteData[127]), .A2(n1193), .B1(
        in_writePathWriteData[127]), .B2(n1188), .ZN(n549) );
  AOI22_X2 U334 ( .A1(in_controlPathWriteData[128]), .A2(n1194), .B1(
        in_writePathWriteData[128]), .B2(n1199), .ZN(n548) );
  AOI22_X2 U336 ( .A1(in_controlPathWriteData[129]), .A2(n1192), .B1(
        in_writePathWriteData[129]), .B2(n1188), .ZN(n547) );
  AOI22_X2 U338 ( .A1(in_controlPathWriteData[130]), .A2(n313), .B1(
        in_writePathWriteData[130]), .B2(n1199), .ZN(n545) );
  AOI22_X2 U340 ( .A1(in_controlPathWriteData[131]), .A2(n1192), .B1(
        in_writePathWriteData[131]), .B2(n1199), .ZN(n544) );
  AOI22_X2 U342 ( .A1(in_controlPathWriteData[132]), .A2(n1193), .B1(
        in_writePathWriteData[132]), .B2(n1199), .ZN(n543) );
  AOI22_X2 U344 ( .A1(in_controlPathWriteData[133]), .A2(n1193), .B1(
        in_writePathWriteData[133]), .B2(n1186), .ZN(n542) );
  AOI22_X2 U346 ( .A1(in_controlPathWriteData[134]), .A2(n313), .B1(
        in_writePathWriteData[134]), .B2(n1186), .ZN(n541) );
  AOI22_X2 U348 ( .A1(in_controlPathWriteData[135]), .A2(n1192), .B1(
        in_writePathWriteData[135]), .B2(n1187), .ZN(n540) );
  AOI22_X2 U350 ( .A1(in_controlPathWriteData[136]), .A2(n1191), .B1(
        in_writePathWriteData[136]), .B2(n1187), .ZN(n539) );
  AOI22_X2 U352 ( .A1(in_controlPathWriteData[137]), .A2(n1193), .B1(
        in_writePathWriteData[137]), .B2(n1186), .ZN(n538) );
  AOI22_X2 U354 ( .A1(in_controlPathWriteData[138]), .A2(n1192), .B1(
        in_writePathWriteData[138]), .B2(n1187), .ZN(n537) );
  AOI22_X2 U356 ( .A1(in_controlPathWriteData[139]), .A2(n1194), .B1(
        in_writePathWriteData[139]), .B2(n1187), .ZN(n536) );
  AOI22_X2 U358 ( .A1(in_controlPathWriteData[140]), .A2(n1193), .B1(
        in_writePathWriteData[140]), .B2(n1189), .ZN(n534) );
  AOI22_X2 U360 ( .A1(in_controlPathWriteData[141]), .A2(n1194), .B1(
        in_writePathWriteData[141]), .B2(n1189), .ZN(n533) );
  AOI22_X2 U362 ( .A1(in_controlPathWriteData[142]), .A2(n1191), .B1(
        in_writePathWriteData[142]), .B2(n1188), .ZN(n532) );
  AOI22_X2 U364 ( .A1(in_controlPathWriteData[143]), .A2(n1194), .B1(
        in_writePathWriteData[143]), .B2(n1186), .ZN(n531) );
  AOI22_X2 U366 ( .A1(in_controlPathWriteData[144]), .A2(n1191), .B1(
        in_writePathWriteData[144]), .B2(n1199), .ZN(n530) );
  AOI22_X2 U368 ( .A1(in_controlPathWriteData[145]), .A2(n1191), .B1(
        in_writePathWriteData[145]), .B2(n1199), .ZN(n529) );
  AOI22_X2 U370 ( .A1(in_controlPathWriteData[146]), .A2(n1194), .B1(
        in_writePathWriteData[146]), .B2(n1189), .ZN(n528) );
  AOI22_X2 U372 ( .A1(in_controlPathWriteData[147]), .A2(n1192), .B1(
        in_writePathWriteData[147]), .B2(n1188), .ZN(n527) );
  AOI22_X2 U374 ( .A1(in_controlPathWriteData[148]), .A2(n1192), .B1(
        in_writePathWriteData[148]), .B2(n1188), .ZN(n526) );
  AOI22_X2 U376 ( .A1(in_controlPathWriteData[149]), .A2(n1192), .B1(
        in_writePathWriteData[149]), .B2(n1186), .ZN(n525) );
  AOI22_X2 U378 ( .A1(in_controlPathWriteData[150]), .A2(n1193), .B1(
        in_writePathWriteData[150]), .B2(n1189), .ZN(n523) );
  AOI22_X2 U380 ( .A1(in_controlPathWriteData[151]), .A2(n1194), .B1(
        in_writePathWriteData[151]), .B2(n1186), .ZN(n522) );
  AOI22_X2 U382 ( .A1(in_controlPathWriteData[152]), .A2(n1191), .B1(
        in_writePathWriteData[152]), .B2(n1188), .ZN(n521) );
  AOI22_X2 U384 ( .A1(in_controlPathWriteData[153]), .A2(n1191), .B1(
        in_writePathWriteData[153]), .B2(n1187), .ZN(n520) );
  AOI22_X2 U386 ( .A1(in_controlPathWriteData[154]), .A2(n1193), .B1(
        in_writePathWriteData[154]), .B2(n1189), .ZN(n519) );
  AOI22_X2 U388 ( .A1(in_controlPathWriteData[155]), .A2(n1192), .B1(
        in_writePathWriteData[155]), .B2(n1187), .ZN(n518) );
  AOI22_X2 U390 ( .A1(in_controlPathWriteData[156]), .A2(n1192), .B1(
        in_writePathWriteData[156]), .B2(n1187), .ZN(n517) );
  AOI22_X2 U392 ( .A1(in_controlPathWriteData[157]), .A2(n1193), .B1(
        in_writePathWriteData[157]), .B2(n1186), .ZN(n516) );
  AOI22_X2 U394 ( .A1(in_controlPathWriteData[158]), .A2(n1194), .B1(
        in_writePathWriteData[158]), .B2(n1188), .ZN(n515) );
  AOI22_X2 U396 ( .A1(in_controlPathWriteData[159]), .A2(n1193), .B1(
        in_writePathWriteData[159]), .B2(n1189), .ZN(n514) );
  AOI22_X2 U398 ( .A1(in_controlPathWriteData[160]), .A2(n1194), .B1(
        in_writePathWriteData[160]), .B2(n1188), .ZN(n512) );
  AOI22_X2 U400 ( .A1(in_controlPathWriteData[161]), .A2(n1193), .B1(
        in_writePathWriteData[161]), .B2(n1189), .ZN(n511) );
  AOI22_X2 U402 ( .A1(in_controlPathWriteData[162]), .A2(n1194), .B1(
        in_writePathWriteData[162]), .B2(n1187), .ZN(n510) );
  AOI22_X2 U404 ( .A1(in_controlPathWriteData[163]), .A2(n1191), .B1(
        in_writePathWriteData[163]), .B2(n1186), .ZN(n509) );
  AOI22_X2 U406 ( .A1(in_controlPathWriteData[164]), .A2(n1194), .B1(
        in_writePathWriteData[164]), .B2(n1188), .ZN(n508) );
  AOI22_X2 U408 ( .A1(in_controlPathWriteData[165]), .A2(n1191), .B1(
        in_writePathWriteData[165]), .B2(n1199), .ZN(n507) );
  AOI22_X2 U410 ( .A1(in_controlPathWriteData[166]), .A2(n1192), .B1(
        in_writePathWriteData[166]), .B2(n1186), .ZN(n506) );
  AOI22_X2 U412 ( .A1(in_controlPathWriteData[167]), .A2(n1191), .B1(
        in_writePathWriteData[167]), .B2(n1199), .ZN(n505) );
  AOI22_X2 U414 ( .A1(in_controlPathWriteData[168]), .A2(n1193), .B1(
        in_writePathWriteData[168]), .B2(n1199), .ZN(n504) );
  AOI22_X2 U416 ( .A1(in_controlPathWriteData[169]), .A2(n1192), .B1(
        in_writePathWriteData[169]), .B2(n1199), .ZN(n503) );
  AOI22_X2 U418 ( .A1(in_controlPathWriteData[170]), .A2(n1192), .B1(
        in_writePathWriteData[170]), .B2(n1199), .ZN(n501) );
  AOI22_X2 U420 ( .A1(in_controlPathWriteData[171]), .A2(n1191), .B1(
        in_writePathWriteData[171]), .B2(n1199), .ZN(n500) );
  AOI22_X2 U422 ( .A1(in_controlPathWriteData[172]), .A2(n1194), .B1(
        in_writePathWriteData[172]), .B2(n1199), .ZN(n499) );
  AOI22_X2 U424 ( .A1(in_controlPathWriteData[173]), .A2(n1192), .B1(
        in_writePathWriteData[173]), .B2(n1199), .ZN(n498) );
  AOI22_X2 U426 ( .A1(in_controlPathWriteData[174]), .A2(n1193), .B1(
        in_writePathWriteData[174]), .B2(n1186), .ZN(n497) );
  AOI22_X2 U428 ( .A1(in_controlPathWriteData[175]), .A2(n1193), .B1(
        in_writePathWriteData[175]), .B2(n1189), .ZN(n496) );
  AOI22_X2 U430 ( .A1(in_controlPathWriteData[176]), .A2(n1194), .B1(
        in_writePathWriteData[176]), .B2(n1187), .ZN(n495) );
  AOI22_X2 U432 ( .A1(in_controlPathWriteData[177]), .A2(n1191), .B1(
        in_writePathWriteData[177]), .B2(n1187), .ZN(n494) );
  AOI22_X2 U434 ( .A1(in_controlPathWriteData[178]), .A2(n1193), .B1(
        in_writePathWriteData[178]), .B2(n1187), .ZN(n493) );
  AOI22_X2 U436 ( .A1(in_controlPathWriteData[179]), .A2(n1194), .B1(
        in_writePathWriteData[179]), .B2(n1189), .ZN(n492) );
  AOI22_X2 U438 ( .A1(in_controlPathWriteData[180]), .A2(n1191), .B1(
        in_writePathWriteData[180]), .B2(n1189), .ZN(n490) );
  AOI22_X2 U440 ( .A1(in_controlPathWriteData[181]), .A2(n1194), .B1(
        in_writePathWriteData[181]), .B2(n1199), .ZN(n489) );
  AOI22_X2 U442 ( .A1(in_controlPathWriteData[182]), .A2(n1191), .B1(
        in_writePathWriteData[182]), .B2(n1188), .ZN(n488) );
  AOI22_X2 U444 ( .A1(in_controlPathWriteData[183]), .A2(n1192), .B1(
        in_writePathWriteData[183]), .B2(n1188), .ZN(n487) );
  AOI22_X2 U446 ( .A1(in_controlPathWriteData[184]), .A2(n1191), .B1(
        in_writePathWriteData[184]), .B2(n1188), .ZN(n486) );
  AOI22_X2 U448 ( .A1(in_controlPathWriteData[185]), .A2(n1192), .B1(
        in_writePathWriteData[185]), .B2(n1189), .ZN(n485) );
  AOI22_X2 U450 ( .A1(in_controlPathWriteData[186]), .A2(n1193), .B1(
        in_writePathWriteData[186]), .B2(n1186), .ZN(n484) );
  AOI22_X2 U452 ( .A1(in_controlPathWriteData[187]), .A2(n1194), .B1(
        in_writePathWriteData[187]), .B2(n1199), .ZN(n483) );
  AOI22_X2 U454 ( .A1(in_controlPathWriteData[188]), .A2(n1192), .B1(
        in_writePathWriteData[188]), .B2(n1188), .ZN(n482) );
  AOI22_X2 U456 ( .A1(in_controlPathWriteData[189]), .A2(n1191), .B1(
        in_writePathWriteData[189]), .B2(n1186), .ZN(n481) );
  AOI22_X2 U458 ( .A1(in_controlPathWriteData[190]), .A2(n1192), .B1(
        in_writePathWriteData[190]), .B2(n1187), .ZN(n479) );
  AOI22_X2 U460 ( .A1(in_controlPathWriteData[191]), .A2(n1193), .B1(
        in_writePathWriteData[191]), .B2(n1186), .ZN(n478) );
  AOI22_X2 U462 ( .A1(in_controlPathWriteData[192]), .A2(n1193), .B1(
        in_writePathWriteData[192]), .B2(n1186), .ZN(n477) );
  AOI22_X2 U464 ( .A1(in_controlPathWriteData[193]), .A2(n1192), .B1(
        in_writePathWriteData[193]), .B2(n1187), .ZN(n476) );
  AOI22_X2 U466 ( .A1(in_controlPathWriteData[194]), .A2(n1193), .B1(
        in_writePathWriteData[194]), .B2(n1187), .ZN(n475) );
  AOI22_X2 U468 ( .A1(in_controlPathWriteData[195]), .A2(n1194), .B1(
        in_writePathWriteData[195]), .B2(n1187), .ZN(n474) );
  AOI22_X2 U470 ( .A1(in_controlPathWriteData[196]), .A2(n1191), .B1(
        in_writePathWriteData[196]), .B2(n1189), .ZN(n473) );
  AOI22_X2 U472 ( .A1(in_controlPathWriteData[197]), .A2(n1193), .B1(
        in_writePathWriteData[197]), .B2(n1189), .ZN(n472) );
  AOI22_X2 U474 ( .A1(in_controlPathWriteData[198]), .A2(n1192), .B1(
        in_writePathWriteData[198]), .B2(n1189), .ZN(n471) );
  AOI22_X2 U476 ( .A1(in_controlPathWriteData[199]), .A2(n1194), .B1(
        in_writePathWriteData[199]), .B2(n1188), .ZN(n470) );
  AOI22_X2 U478 ( .A1(in_controlPathWriteData[200]), .A2(n1191), .B1(
        in_writePathWriteData[200]), .B2(n1189), .ZN(n467) );
  AOI22_X2 U480 ( .A1(in_controlPathWriteData[201]), .A2(n1194), .B1(
        in_writePathWriteData[201]), .B2(n1188), .ZN(n466) );
  AOI22_X2 U482 ( .A1(in_controlPathWriteData[202]), .A2(n1194), .B1(
        in_writePathWriteData[202]), .B2(n1188), .ZN(n465) );
  AOI22_X2 U484 ( .A1(in_controlPathWriteData[203]), .A2(n1192), .B1(
        in_writePathWriteData[203]), .B2(n1199), .ZN(n464) );
  AOI22_X2 U486 ( .A1(in_controlPathWriteData[204]), .A2(n1193), .B1(
        in_writePathWriteData[204]), .B2(n1186), .ZN(n463) );
  AOI22_X2 U488 ( .A1(in_controlPathWriteData[205]), .A2(n1194), .B1(
        in_writePathWriteData[205]), .B2(n1199), .ZN(n462) );
  AOI22_X2 U490 ( .A1(in_controlPathWriteData[206]), .A2(n1191), .B1(
        in_writePathWriteData[206]), .B2(n1186), .ZN(n461) );
  AOI22_X2 U492 ( .A1(in_controlPathWriteData[207]), .A2(n1191), .B1(
        in_writePathWriteData[207]), .B2(n1187), .ZN(n460) );
  AOI22_X2 U494 ( .A1(in_controlPathWriteData[208]), .A2(n1193), .B1(
        in_writePathWriteData[208]), .B2(n1189), .ZN(n459) );
  AOI22_X2 U496 ( .A1(in_controlPathWriteData[209]), .A2(n1194), .B1(
        in_writePathWriteData[209]), .B2(n1188), .ZN(n458) );
  AOI22_X2 U498 ( .A1(in_controlPathWriteData[210]), .A2(n1192), .B1(
        in_writePathWriteData[210]), .B2(n1186), .ZN(n456) );
  AOI22_X2 U500 ( .A1(in_controlPathWriteData[211]), .A2(n1191), .B1(
        in_writePathWriteData[211]), .B2(n1187), .ZN(n455) );
  AOI22_X2 U502 ( .A1(in_controlPathWriteData[212]), .A2(n1192), .B1(
        in_writePathWriteData[212]), .B2(n1189), .ZN(n454) );
  AOI22_X2 U504 ( .A1(in_controlPathWriteData[213]), .A2(n313), .B1(
        in_writePathWriteData[213]), .B2(n1188), .ZN(n453) );
  AOI22_X2 U506 ( .A1(in_controlPathWriteData[214]), .A2(n1191), .B1(
        in_writePathWriteData[214]), .B2(n1186), .ZN(n452) );
  AOI22_X2 U508 ( .A1(in_controlPathWriteData[215]), .A2(n313), .B1(
        in_writePathWriteData[215]), .B2(n1187), .ZN(n451) );
  AOI22_X2 U510 ( .A1(in_controlPathWriteData[216]), .A2(n1192), .B1(
        in_writePathWriteData[216]), .B2(n1189), .ZN(n450) );
  AOI22_X2 U512 ( .A1(in_controlPathWriteData[217]), .A2(n1193), .B1(
        in_writePathWriteData[217]), .B2(n1188), .ZN(n449) );
  AOI22_X2 U514 ( .A1(in_controlPathWriteData[218]), .A2(n1193), .B1(
        in_writePathWriteData[218]), .B2(n1186), .ZN(n448) );
  AOI22_X2 U516 ( .A1(in_controlPathWriteData[219]), .A2(n1194), .B1(
        in_writePathWriteData[219]), .B2(n1187), .ZN(n447) );
  AOI22_X2 U518 ( .A1(in_controlPathWriteData[220]), .A2(n1193), .B1(
        in_writePathWriteData[220]), .B2(n1189), .ZN(n445) );
  AOI22_X2 U520 ( .A1(in_controlPathWriteData[221]), .A2(n1192), .B1(
        in_writePathWriteData[221]), .B2(n1188), .ZN(n444) );
  AOI22_X2 U522 ( .A1(in_controlPathWriteData[222]), .A2(n313), .B1(
        in_writePathWriteData[222]), .B2(n1186), .ZN(n443) );
  AOI22_X2 U524 ( .A1(in_controlPathWriteData[223]), .A2(n1194), .B1(
        in_writePathWriteData[223]), .B2(n1187), .ZN(n442) );
  AOI22_X2 U526 ( .A1(in_controlPathWriteData[224]), .A2(n1191), .B1(
        in_writePathWriteData[224]), .B2(n1189), .ZN(n441) );
  AOI22_X2 U528 ( .A1(in_controlPathWriteData[225]), .A2(n1192), .B1(
        in_writePathWriteData[225]), .B2(n1188), .ZN(n440) );
  AOI22_X2 U530 ( .A1(in_controlPathWriteData[226]), .A2(n1191), .B1(
        in_writePathWriteData[226]), .B2(n1186), .ZN(n439) );
  AOI22_X2 U532 ( .A1(in_controlPathWriteData[227]), .A2(n1192), .B1(
        in_writePathWriteData[227]), .B2(n1187), .ZN(n438) );
  AOI22_X2 U534 ( .A1(in_controlPathWriteData[228]), .A2(n1193), .B1(
        in_writePathWriteData[228]), .B2(n1188), .ZN(n437) );
  AOI22_X2 U536 ( .A1(in_controlPathWriteData[229]), .A2(n1193), .B1(
        in_writePathWriteData[229]), .B2(n1186), .ZN(n436) );
  AOI22_X2 U538 ( .A1(in_controlPathWriteData[230]), .A2(n1194), .B1(
        in_writePathWriteData[230]), .B2(n1187), .ZN(n434) );
  AOI22_X2 U540 ( .A1(in_controlPathWriteData[231]), .A2(n1194), .B1(
        in_writePathWriteData[231]), .B2(n1189), .ZN(n433) );
  AOI22_X2 U542 ( .A1(in_controlPathWriteData[232]), .A2(n1191), .B1(
        in_writePathWriteData[232]), .B2(n1186), .ZN(n432) );
  AOI22_X2 U544 ( .A1(in_controlPathWriteData[233]), .A2(n313), .B1(
        in_writePathWriteData[233]), .B2(n1187), .ZN(n431) );
  AOI22_X2 U546 ( .A1(in_controlPathWriteData[234]), .A2(n1194), .B1(
        in_writePathWriteData[234]), .B2(n1189), .ZN(n430) );
  AOI22_X2 U548 ( .A1(in_controlPathWriteData[235]), .A2(n1193), .B1(
        in_writePathWriteData[235]), .B2(n1188), .ZN(n429) );
  AOI22_X2 U550 ( .A1(in_controlPathWriteData[236]), .A2(n1191), .B1(
        in_writePathWriteData[236]), .B2(n1187), .ZN(n428) );
  AOI22_X2 U552 ( .A1(in_controlPathWriteData[237]), .A2(n313), .B1(
        in_writePathWriteData[237]), .B2(n1189), .ZN(n427) );
  AOI22_X2 U554 ( .A1(in_controlPathWriteData[238]), .A2(n313), .B1(
        in_writePathWriteData[238]), .B2(n1188), .ZN(n426) );
  AOI22_X2 U556 ( .A1(in_controlPathWriteData[239]), .A2(n1192), .B1(
        in_writePathWriteData[239]), .B2(n1188), .ZN(n425) );
  AOI22_X2 U558 ( .A1(in_controlPathWriteData[240]), .A2(n1191), .B1(
        in_writePathWriteData[240]), .B2(n1186), .ZN(n423) );
  AOI22_X2 U560 ( .A1(in_controlPathWriteData[241]), .A2(n1194), .B1(
        in_writePathWriteData[241]), .B2(n1187), .ZN(n422) );
  AOI22_X2 U562 ( .A1(in_controlPathWriteData[242]), .A2(n1191), .B1(
        in_writePathWriteData[242]), .B2(n1189), .ZN(n421) );
  AOI22_X2 U564 ( .A1(in_controlPathWriteData[243]), .A2(n1192), .B1(
        in_writePathWriteData[243]), .B2(n1188), .ZN(n420) );
  AOI22_X2 U566 ( .A1(in_controlPathWriteData[244]), .A2(n1192), .B1(
        in_writePathWriteData[244]), .B2(n1186), .ZN(n419) );
  AOI22_X2 U568 ( .A1(in_controlPathWriteData[245]), .A2(n313), .B1(
        in_writePathWriteData[245]), .B2(n1187), .ZN(n418) );
  AOI22_X2 U570 ( .A1(in_controlPathWriteData[246]), .A2(n313), .B1(
        in_writePathWriteData[246]), .B2(n1189), .ZN(n417) );
  AOI22_X2 U572 ( .A1(in_controlPathWriteData[247]), .A2(n1193), .B1(
        in_writePathWriteData[247]), .B2(n1188), .ZN(n416) );
  AOI22_X2 U574 ( .A1(in_controlPathWriteData[248]), .A2(n1192), .B1(
        in_writePathWriteData[248]), .B2(n1186), .ZN(n415) );
  AOI22_X2 U576 ( .A1(in_controlPathWriteData[249]), .A2(n1193), .B1(
        in_writePathWriteData[249]), .B2(n1187), .ZN(n414) );
  AOI22_X2 U578 ( .A1(in_controlPathWriteData[250]), .A2(n1194), .B1(
        in_writePathWriteData[250]), .B2(n1199), .ZN(n412) );
  AOI22_X2 U580 ( .A1(in_controlPathWriteData[251]), .A2(n1194), .B1(
        in_writePathWriteData[251]), .B2(n1199), .ZN(n411) );
  AOI22_X2 U582 ( .A1(in_controlPathWriteData[252]), .A2(n1193), .B1(
        in_writePathWriteData[252]), .B2(n1199), .ZN(n410) );
  AOI22_X2 U584 ( .A1(in_controlPathWriteData[253]), .A2(n1191), .B1(
        in_writePathWriteData[253]), .B2(n1199), .ZN(n409) );
  AOI22_X2 U585 ( .A1(in_controlPathWriteData[254]), .A2(n1193), .B1(
        in_writePathWriteData[254]), .B2(n1199), .ZN(n408) );
  AOI22_X2 U588 ( .A1(in_controlPathWriteData[255]), .A2(n1191), .B1(
        in_writePathWriteData[255]), .B2(n1199), .ZN(n407) );
  AOI22_X2 U589 ( .A1(in_controlPathWE), .A2(n313), .B1(in_writePathWE), .B2(
        n1189), .ZN(n312) );
  AOI22_X2 U590 ( .A1(in_controlPathWriteData[96]), .A2(n313), .B1(
        in_writePathWriteData[96]), .B2(n1189), .ZN(n329) );
  AOI22_X2 U591 ( .A1(in_controlPathWriteData[97]), .A2(n313), .B1(
        in_writePathWriteData[97]), .B2(n1186), .ZN(n328) );
  AOI22_X2 U592 ( .A1(in_controlPathWriteData[98]), .A2(n313), .B1(
        in_writePathWriteData[98]), .B2(n1188), .ZN(n327) );
  AOI22_X2 U593 ( .A1(in_controlPathWriteData[99]), .A2(n313), .B1(
        in_writePathWriteData[99]), .B2(n1188), .ZN(n326) );
  AOI22_X2 U594 ( .A1(in_controlPathReadAddr2[0]), .A2(n1184), .B1(
        in_writePathReadAddr2[0]), .B2(n1185), .ZN(n310) );
  AOI22_X2 U595 ( .A1(in_controlPathReadAddr2[3]), .A2(n1184), .B1(
        in_writePathReadAddr2[3]), .B2(n1185), .ZN(n306) );
  AOI22_X2 U596 ( .A1(in_controlPathReadAddr2[5]), .A2(n1184), .B1(
        in_writePathReadAddr2[5]), .B2(n1185), .ZN(n304) );
  AOI22_X2 U597 ( .A1(in_controlPathReadAddr2[7]), .A2(n1184), .B1(
        in_writePathReadAddr2[7]), .B2(n1185), .ZN(n302) );
  AOI22_X2 U598 ( .A1(in_controlPathReadAddr2[8]), .A2(n1184), .B1(
        in_writePathReadAddr2[8]), .B2(n1185), .ZN(n301) );
  AOI22_X2 U599 ( .A1(in_controlPathReadAddr2[9]), .A2(n1184), .B1(
        in_writePathReadAddr2[9]), .B2(n1185), .ZN(n299) );
  AOI22_X2 U600 ( .A1(in_controlPathReadAddr2[10]), .A2(n1184), .B1(
        in_writePathReadAddr2[10]), .B2(n1185), .ZN(n308) );
  INV_X4 U601 ( .A(n288), .ZN(n1197) );
  OAI211_X2 U602 ( .C1(in_yWriteModuleEnable), .C2(in_yComputeModuleEnable), 
        .A(n311), .B(reset), .ZN(n288) );
  INV_X8 U38 ( .A(n1190), .ZN(n1188) );
  INV_X8 U42 ( .A(n1190), .ZN(n1189) );
  INV_X8 U46 ( .A(n1190), .ZN(n1187) );
  INV_X8 U48 ( .A(n1190), .ZN(n1186) );
  INV_X1 U71 ( .A(n1183), .ZN(n1198) );
  INV_X8 U74 ( .A(n1198), .ZN(n1199) );
  INV_X8 U76 ( .A(n1195), .ZN(n1191) );
  INV_X8 U78 ( .A(n1195), .ZN(n1194) );
  INV_X8 U603 ( .A(n1195), .ZN(n1193) );
  INV_X8 U604 ( .A(n1195), .ZN(n1192) );
endmodule


module busWriteY ( clock, reset, inModuleEnable, cpDoneFlag, dpDoneFlag, 
        inDiagAddr, inNonDAddr, inDiagOH, inNonDiagOH, inYreadData1, 
        inYreadData2, inYComputedVal, inYchngData, op_writeData, 
        op_writeAddress, op_readStoreAddr, op_WEbit, op_writeDone );
  input [10:0] inDiagAddr;
  input [10:0] inNonDAddr;
  input [3:0] inDiagOH;
  input [3:0] inNonDiagOH;
  input [255:0] inYreadData1;
  input [255:0] inYreadData2;
  input [47:0] inYComputedVal;
  input [47:0] inYchngData;
  output [255:0] op_writeData;
  output [10:0] op_writeAddress;
  output [10:0] op_readStoreAddr;
  input clock, reset, inModuleEnable, cpDoneFlag, dpDoneFlag;
  output op_WEbit, op_writeDone;
  wire   n1799, U62_Z_0, U62_Z_1, U62_Z_2, U62_Z_3, U62_Z_4, U62_Z_5, U62_Z_6,
         U62_Z_7, U62_Z_8, U62_Z_9, U62_Z_10, U62_Z_11, U62_Z_12, U62_Z_13,
         U62_Z_14, U62_Z_15, U62_Z_16, U62_Z_17, U62_Z_18, U62_Z_19, U62_Z_20,
         U62_Z_21, U62_Z_22, U62_Z_23, U62_Z_24, U62_Z_25, U62_Z_26, U62_Z_27,
         U62_Z_28, U62_Z_29, U62_Z_30, U62_Z_31, U62_Z_32, U62_Z_33, U62_Z_34,
         U62_Z_35, U62_Z_36, U62_Z_37, U62_Z_38, U62_Z_39, U62_Z_40, U62_Z_41,
         U62_Z_42, U62_Z_43, U62_Z_44, U62_Z_45, U62_Z_46, U62_Z_47, U62_Z_64,
         U62_Z_65, U62_Z_66, U62_Z_67, U62_Z_68, U62_Z_69, U62_Z_70, U62_Z_71,
         U62_Z_72, U62_Z_73, U62_Z_74, U62_Z_75, U62_Z_76, U62_Z_77, U62_Z_78,
         U62_Z_79, U62_Z_80, U62_Z_81, U62_Z_82, U62_Z_83, U62_Z_84, U62_Z_85,
         U62_Z_86, U62_Z_87, U62_Z_88, U62_Z_89, U62_Z_90, U62_Z_91, U62_Z_92,
         U62_Z_93, U62_Z_94, U62_Z_95, U62_Z_96, U62_Z_97, U62_Z_98, U62_Z_99,
         U62_Z_100, U62_Z_101, U62_Z_102, U62_Z_103, U62_Z_104, U62_Z_105,
         U62_Z_106, U62_Z_107, U62_Z_108, U62_Z_109, U62_Z_110, U62_Z_111,
         U62_Z_128, U62_Z_129, U62_Z_130, U62_Z_131, U62_Z_132, U62_Z_133,
         U62_Z_134, U62_Z_135, U62_Z_136, U62_Z_137, U62_Z_138, U62_Z_139,
         U62_Z_140, U62_Z_141, U62_Z_142, U62_Z_143, U62_Z_144, U62_Z_145,
         U62_Z_146, U62_Z_147, U62_Z_148, U62_Z_149, U62_Z_150, U62_Z_151,
         U62_Z_152, U62_Z_153, U62_Z_154, U62_Z_155, U62_Z_156, U62_Z_157,
         U62_Z_158, U62_Z_159, U62_Z_160, U62_Z_161, U62_Z_162, U62_Z_163,
         U62_Z_164, U62_Z_165, U62_Z_166, U62_Z_167, U62_Z_168, U62_Z_169,
         U62_Z_170, U62_Z_171, U62_Z_172, U62_Z_173, U62_Z_174, U62_Z_175,
         U61_Z_0, U61_Z_1, U61_Z_2, U61_Z_3, U61_Z_4, U61_Z_5, U61_Z_6,
         U61_Z_7, U61_Z_8, U61_Z_9, U61_Z_10, U59_Z_0, U59_Z_1, U59_Z_2,
         U59_Z_3, U59_Z_4, U59_Z_5, U59_Z_6, U59_Z_7, U59_Z_8, U59_Z_9,
         U59_Z_10, U58_Z_0, U57_Z_0, U57_Z_1, U57_Z_2, U57_Z_3, U57_Z_4,
         U57_Z_5, U57_Z_6, U57_Z_7, U57_Z_8, U57_Z_9, U57_Z_10, U57_Z_11,
         U57_Z_12, U57_Z_13, U57_Z_14, U57_Z_15, U57_Z_16, U57_Z_17, U57_Z_18,
         U57_Z_19, U57_Z_20, U57_Z_21, U57_Z_22, U57_Z_23, U57_Z_24, U57_Z_25,
         U57_Z_26, U57_Z_27, U57_Z_28, U57_Z_29, U57_Z_30, U57_Z_31, U57_Z_32,
         U57_Z_33, U57_Z_34, U57_Z_35, U57_Z_36, U57_Z_37, U57_Z_38, U57_Z_39,
         U57_Z_40, U57_Z_41, U57_Z_42, U57_Z_43, U57_Z_44, U57_Z_45, U57_Z_46,
         U57_Z_47, U57_Z_48, U57_Z_49, U57_Z_50, U57_Z_51, U57_Z_52, U57_Z_53,
         U57_Z_54, U57_Z_55, U57_Z_56, U57_Z_57, U57_Z_58, U57_Z_59, U57_Z_60,
         U57_Z_61, U57_Z_62, U57_Z_63, U57_Z_64, U57_Z_65, U57_Z_66, U57_Z_67,
         U57_Z_68, U57_Z_69, U57_Z_70, U57_Z_71, U57_Z_72, U57_Z_73, U57_Z_74,
         U57_Z_75, U57_Z_76, U57_Z_77, U57_Z_78, U57_Z_79, U57_Z_80, U57_Z_81,
         U57_Z_82, U57_Z_83, U57_Z_84, U57_Z_85, U57_Z_86, U57_Z_87, U57_Z_88,
         U57_Z_89, U57_Z_90, U57_Z_91, U57_Z_92, U57_Z_93, U57_Z_94, U57_Z_95,
         U57_Z_96, U57_Z_97, U57_Z_98, U57_Z_99, U57_Z_100, U57_Z_101,
         U57_Z_102, U57_Z_103, U57_Z_104, U57_Z_105, U57_Z_106, U57_Z_107,
         U57_Z_108, U57_Z_109, U57_Z_110, U57_Z_111, U57_Z_112, U57_Z_113,
         U57_Z_114, U57_Z_115, U57_Z_116, U57_Z_117, U57_Z_118, U57_Z_119,
         U57_Z_120, U57_Z_121, U57_Z_122, U57_Z_123, U57_Z_124, U57_Z_125,
         U57_Z_126, U57_Z_127, U57_Z_128, U57_Z_129, U57_Z_130, U57_Z_131,
         U57_Z_132, U57_Z_133, U57_Z_134, U57_Z_135, U57_Z_136, U57_Z_137,
         U57_Z_138, U57_Z_139, U57_Z_140, U57_Z_141, U57_Z_142, U57_Z_143,
         U57_Z_144, U57_Z_145, U57_Z_146, U57_Z_147, U57_Z_148, U57_Z_149,
         U57_Z_150, U57_Z_151, U57_Z_152, U57_Z_153, U57_Z_154, U57_Z_155,
         U57_Z_156, U57_Z_157, U57_Z_158, U57_Z_159, U57_Z_160, U57_Z_161,
         U57_Z_162, U57_Z_163, U57_Z_164, U57_Z_165, U57_Z_166, U57_Z_167,
         U57_Z_168, U57_Z_169, U57_Z_170, U57_Z_171, U57_Z_172, U57_Z_173,
         U57_Z_174, U57_Z_175, U57_Z_176, U57_Z_177, U57_Z_178, U57_Z_179,
         U57_Z_180, U57_Z_181, U57_Z_182, U57_Z_183, U57_Z_184, U57_Z_185,
         U57_Z_186, U57_Z_187, U57_Z_188, U57_Z_189, U57_Z_190, U57_Z_191,
         U57_Z_192, U57_Z_193, U57_Z_194, U57_Z_195, U57_Z_196, U57_Z_197,
         U57_Z_198, U57_Z_199, U57_Z_200, U57_Z_201, U57_Z_202, U57_Z_203,
         U57_Z_204, U57_Z_205, U57_Z_206, U57_Z_207, U57_Z_208, U57_Z_209,
         U57_Z_210, U57_Z_211, U57_Z_212, U57_Z_213, U57_Z_214, U57_Z_215,
         U57_Z_216, U57_Z_217, U57_Z_218, U57_Z_219, U57_Z_220, U57_Z_221,
         U57_Z_222, U57_Z_223, U57_Z_224, U57_Z_225, U57_Z_226, U57_Z_227,
         U57_Z_228, U57_Z_229, U57_Z_230, U57_Z_231, U57_Z_232, U57_Z_233,
         U57_Z_234, U57_Z_235, U57_Z_236, U57_Z_237, U57_Z_238, U57_Z_239,
         U57_Z_240, U57_Z_241, U57_Z_242, U57_Z_243, U57_Z_244, U57_Z_245,
         U57_Z_246, U57_Z_247, U57_Z_248, U57_Z_249, U57_Z_250, U57_Z_251,
         U57_Z_252, U57_Z_253, U57_Z_254, U57_Z_255, U55_Z_0, U55_Z_1,
         U41_DATA2_0, U41_DATA2_1, U41_DATA2_2, U41_DATA2_3, U41_DATA2_4,
         U41_DATA2_5, U41_DATA2_6, U41_DATA2_7, U41_DATA2_8, U41_DATA2_9,
         U41_DATA2_10, U41_DATA1_0, U41_DATA1_1, U41_DATA1_2, U41_DATA1_3,
         U41_DATA1_4, U41_DATA1_5, U41_DATA1_6, U41_DATA1_7, U41_DATA1_8,
         U41_DATA1_9, U41_DATA1_10, U36_DATA2_0, U36_DATA2_1, U36_DATA2_2,
         U36_DATA2_3, U36_DATA1_0, U36_DATA1_1, U36_DATA1_2, U36_DATA1_3,
         U35_DATA2_0, U35_DATA2_1, U35_DATA2_2, U35_DATA2_3, U35_DATA1_0,
         U35_DATA1_1, U35_DATA1_2, U35_DATA1_3, U6_DATA3_48, U6_DATA3_49,
         U6_DATA3_50, U6_DATA3_51, U6_DATA3_52, U6_DATA3_53, U6_DATA3_54,
         U6_DATA3_55, U6_DATA3_56, U6_DATA3_57, U6_DATA3_58, U6_DATA3_59,
         U6_DATA3_60, U6_DATA3_61, U6_DATA3_62, U6_DATA3_63, U6_DATA3_112,
         U6_DATA3_113, U6_DATA3_114, U6_DATA3_115, U6_DATA3_116, U6_DATA3_117,
         U6_DATA3_118, U6_DATA3_119, U6_DATA3_120, U6_DATA3_121, U6_DATA3_122,
         U6_DATA3_123, U6_DATA3_124, U6_DATA3_125, U6_DATA3_126, U6_DATA3_127,
         U6_DATA3_176, U6_DATA3_177, U6_DATA3_178, U6_DATA3_179, U6_DATA3_180,
         U6_DATA3_181, U6_DATA3_182, U6_DATA3_183, U6_DATA3_184, U6_DATA3_185,
         U6_DATA3_186, U6_DATA3_187, U6_DATA3_188, U6_DATA3_189, U6_DATA3_190,
         U6_DATA3_191, U6_DATA3_192, U6_DATA3_193, U6_DATA3_194, U6_DATA3_195,
         U6_DATA3_196, U6_DATA3_197, U6_DATA3_198, U6_DATA3_199, U6_DATA3_200,
         U6_DATA3_201, U6_DATA3_202, U6_DATA3_203, U6_DATA3_204, U6_DATA3_205,
         U6_DATA3_206, U6_DATA3_207, U6_DATA3_208, U6_DATA3_209, U6_DATA3_210,
         U6_DATA3_211, U6_DATA3_212, U6_DATA3_213, U6_DATA3_214, U6_DATA3_215,
         U6_DATA3_216, U6_DATA3_217, U6_DATA3_218, U6_DATA3_219, U6_DATA3_220,
         U6_DATA3_221, U6_DATA3_222, U6_DATA3_223, U6_DATA3_224, U6_DATA3_225,
         U6_DATA3_226, U6_DATA3_227, U6_DATA3_228, U6_DATA3_229, U6_DATA3_230,
         U6_DATA3_231, U6_DATA3_232, U6_DATA3_233, U6_DATA3_234, U6_DATA3_235,
         U6_DATA3_236, U6_DATA3_237, U6_DATA3_238, U6_DATA3_239, U6_DATA3_240,
         U6_DATA3_241, U6_DATA3_242, U6_DATA3_243, U6_DATA3_244, U6_DATA3_245,
         U6_DATA3_246, U6_DATA3_247, U6_DATA3_248, U6_DATA3_249, U6_DATA3_250,
         U6_DATA3_251, U6_DATA3_252, U6_DATA3_253, U6_DATA3_254, U6_DATA3_255,
         n4, n5, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n780,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1187, n1190, n1191, n1192, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333;
  wire   [3037:3036] n;

  SDFF_X1 tempDPFlag_reg ( .D(dpDoneFlag), .SI(1'b0), .SE(n4321), .CK(clock), 
        .QN(n4) );
  SDFF_X1 tempCPFlag_reg ( .D(cpDoneFlag), .SI(1'b0), .SE(n4321), .CK(clock), 
        .Q(n1799) );
  DFF_X1 current_state_reg_0_ ( .D(U55_Z_0), .CK(clock), .Q(n[3036]) );
  DFF_X2 tempDiagAddr1_reg_0_ ( .D(n1372), .CK(clock), .QN(n297) );
  DFF_X2 tempDiagAddr1_reg_1_ ( .D(n1373), .CK(clock), .QN(n296) );
  DFF_X2 tempDiagAddr1_reg_2_ ( .D(n1374), .CK(clock), .QN(n295) );
  DFF_X2 tempDiagAddr1_reg_3_ ( .D(n1375), .CK(clock), .QN(n294) );
  DFF_X2 tempDiagAddr1_reg_4_ ( .D(n1376), .CK(clock), .QN(n293) );
  DFF_X2 tempDiagAddr1_reg_5_ ( .D(n1377), .CK(clock), .QN(n292) );
  DFF_X2 tempDiagAddr1_reg_6_ ( .D(n1378), .CK(clock), .QN(n291) );
  DFF_X2 tempDiagAddr1_reg_7_ ( .D(n1379), .CK(clock), .QN(n290) );
  DFF_X2 tempDiagAddr1_reg_8_ ( .D(n1380), .CK(clock), .QN(n289) );
  DFF_X2 tempDiagAddr1_reg_9_ ( .D(n1381), .CK(clock), .QN(n288) );
  DFF_X2 tempDiagAddr1_reg_10_ ( .D(n1382), .CK(clock), .QN(n287) );
  DFF_X2 tempDiagAddr2_reg_0_ ( .D(n1350), .CK(clock), .QN(n308) );
  DFF_X2 tempDiagAddr2_reg_1_ ( .D(n1351), .CK(clock), .QN(n307) );
  DFF_X2 tempDiagAddr2_reg_2_ ( .D(n1352), .CK(clock), .QN(n306) );
  DFF_X2 tempDiagAddr2_reg_3_ ( .D(n1353), .CK(clock), .QN(n305) );
  DFF_X2 tempDiagAddr2_reg_4_ ( .D(n1354), .CK(clock), .QN(n304) );
  DFF_X2 tempDiagAddr2_reg_5_ ( .D(n1355), .CK(clock), .QN(n303) );
  DFF_X2 tempDiagAddr2_reg_6_ ( .D(n1356), .CK(clock), .QN(n302) );
  DFF_X2 tempDiagAddr2_reg_7_ ( .D(n1357), .CK(clock), .QN(n301) );
  DFF_X2 tempDiagAddr2_reg_8_ ( .D(n1358), .CK(clock), .QN(n300) );
  DFF_X2 tempDiagAddr2_reg_9_ ( .D(n1359), .CK(clock), .QN(n299) );
  DFF_X2 tempDiagAddr2_reg_10_ ( .D(n1360), .CK(clock), .QN(n298) );
  DFF_X1 op_readStoreAddr_reg_0_ ( .D(U59_Z_0), .CK(clock), .Q(
        op_readStoreAddr[0]) );
  SDFF_X1 op_WEbit_reg ( .D(n[3037]), .SI(1'b0), .SE(n4290), .CK(clock), .Q(
        op_WEbit) );
  DFF_X1 op_readStoreAddr_reg_3_ ( .D(U59_Z_3), .CK(clock), .Q(
        op_readStoreAddr[3]) );
  DFF_X1 op_writeAddress_reg_3_ ( .D(U61_Z_3), .CK(clock), .Q(
        op_writeAddress[3]) );
  DFF_X1 op_readStoreAddr_reg_5_ ( .D(U59_Z_5), .CK(clock), .Q(
        op_readStoreAddr[5]) );
  DFF_X1 op_writeAddress_reg_5_ ( .D(U61_Z_5), .CK(clock), .Q(
        op_writeAddress[5]) );
  DFF_X1 op_readStoreAddr_reg_4_ ( .D(U59_Z_4), .CK(clock), .Q(
        op_readStoreAddr[4]) );
  DFF_X1 op_writeAddress_reg_4_ ( .D(U61_Z_4), .CK(clock), .Q(
        op_writeAddress[4]) );
  DFF_X1 op_readStoreAddr_reg_1_ ( .D(U59_Z_1), .CK(clock), .Q(
        op_readStoreAddr[1]) );
  DFF_X1 op_writeAddress_reg_1_ ( .D(U61_Z_1), .CK(clock), .Q(
        op_writeAddress[1]) );
  DFF_X1 op_readStoreAddr_reg_2_ ( .D(U59_Z_2), .CK(clock), .Q(
        op_readStoreAddr[2]) );
  DFF_X1 op_writeAddress_reg_2_ ( .D(U61_Z_2), .CK(clock), .Q(
        op_writeAddress[2]) );
  DFF_X1 op_readStoreAddr_reg_6_ ( .D(U59_Z_6), .CK(clock), .Q(
        op_readStoreAddr[6]) );
  DFF_X1 op_writeAddress_reg_6_ ( .D(U61_Z_6), .CK(clock), .Q(
        op_writeAddress[6]) );
  DFF_X1 op_readStoreAddr_reg_8_ ( .D(U59_Z_8), .CK(clock), .Q(
        op_readStoreAddr[8]) );
  DFF_X1 op_writeAddress_reg_8_ ( .D(U61_Z_8), .CK(clock), .Q(
        op_writeAddress[8]) );
  DFF_X1 op_writeAddress_reg_7_ ( .D(U61_Z_7), .CK(clock), .Q(
        op_writeAddress[7]) );
  DFF_X1 op_readStoreAddr_reg_7_ ( .D(U59_Z_7), .CK(clock), .Q(
        op_readStoreAddr[7]) );
  DFF_X1 op_readStoreAddr_reg_9_ ( .D(U59_Z_9), .CK(clock), .Q(
        op_readStoreAddr[9]) );
  DFF_X1 op_writeAddress_reg_9_ ( .D(U61_Z_9), .CK(clock), .Q(
        op_writeAddress[9]) );
  DFF_X1 op_readStoreAddr_reg_10_ ( .D(U59_Z_10), .CK(clock), .Q(
        op_readStoreAddr[10]) );
  DFF_X1 op_writeAddress_reg_10_ ( .D(U61_Z_10), .CK(clock), .Q(
        op_writeAddress[10]) );
  DFF_X1 op_writeDone_reg ( .D(U58_Z_0), .CK(clock), .Q(op_writeDone) );
  DFF_X1 op_writeAddress_reg_0_ ( .D(U61_Z_0), .CK(clock), .Q(
        op_writeAddress[0]) );
  DFF_X1 tempStoreData_reg_239_ ( .D(U57_Z_239), .CK(clock), .Q(U6_DATA3_239)
         );
  DFF_X1 tempStoreData_reg_238_ ( .D(U57_Z_238), .CK(clock), .Q(U6_DATA3_238)
         );
  DFF_X1 tempStoreData_reg_237_ ( .D(U57_Z_237), .CK(clock), .Q(U6_DATA3_237)
         );
  DFF_X1 tempStoreData_reg_236_ ( .D(U57_Z_236), .CK(clock), .Q(U6_DATA3_236)
         );
  DFF_X1 tempStoreData_reg_235_ ( .D(U57_Z_235), .CK(clock), .Q(U6_DATA3_235)
         );
  DFF_X1 tempStoreData_reg_234_ ( .D(U57_Z_234), .CK(clock), .Q(U6_DATA3_234)
         );
  DFF_X1 tempStoreData_reg_233_ ( .D(U57_Z_233), .CK(clock), .Q(U6_DATA3_233)
         );
  DFF_X1 tempStoreData_reg_232_ ( .D(U57_Z_232), .CK(clock), .Q(U6_DATA3_232)
         );
  DFF_X1 tempStoreData_reg_231_ ( .D(U57_Z_231), .CK(clock), .Q(U6_DATA3_231)
         );
  DFF_X1 tempStoreData_reg_230_ ( .D(U57_Z_230), .CK(clock), .Q(U6_DATA3_230)
         );
  DFF_X1 tempStoreData_reg_229_ ( .D(U57_Z_229), .CK(clock), .Q(U6_DATA3_229)
         );
  DFF_X1 tempStoreData_reg_228_ ( .D(U57_Z_228), .CK(clock), .Q(U6_DATA3_228)
         );
  DFF_X1 tempStoreData_reg_227_ ( .D(U57_Z_227), .CK(clock), .Q(U6_DATA3_227)
         );
  DFF_X1 tempStoreData_reg_226_ ( .D(U57_Z_226), .CK(clock), .Q(U6_DATA3_226)
         );
  DFF_X1 tempStoreData_reg_225_ ( .D(U57_Z_225), .CK(clock), .Q(U6_DATA3_225)
         );
  DFF_X1 tempStoreData_reg_224_ ( .D(U57_Z_224), .CK(clock), .Q(U6_DATA3_224)
         );
  DFF_X1 tempStoreData_reg_223_ ( .D(U57_Z_223), .CK(clock), .Q(U6_DATA3_223)
         );
  DFF_X1 tempStoreData_reg_222_ ( .D(U57_Z_222), .CK(clock), .Q(U6_DATA3_222)
         );
  DFF_X1 tempStoreData_reg_221_ ( .D(U57_Z_221), .CK(clock), .Q(U6_DATA3_221)
         );
  DFF_X1 tempStoreData_reg_220_ ( .D(U57_Z_220), .CK(clock), .Q(U6_DATA3_220)
         );
  DFF_X1 tempStoreData_reg_219_ ( .D(U57_Z_219), .CK(clock), .Q(U6_DATA3_219)
         );
  DFF_X1 tempStoreData_reg_218_ ( .D(U57_Z_218), .CK(clock), .Q(U6_DATA3_218)
         );
  DFF_X1 tempStoreData_reg_217_ ( .D(U57_Z_217), .CK(clock), .Q(U6_DATA3_217)
         );
  DFF_X1 tempStoreData_reg_216_ ( .D(U57_Z_216), .CK(clock), .Q(U6_DATA3_216)
         );
  DFF_X1 tempStoreData_reg_215_ ( .D(U57_Z_215), .CK(clock), .Q(U6_DATA3_215)
         );
  DFF_X1 tempStoreData_reg_214_ ( .D(U57_Z_214), .CK(clock), .Q(U6_DATA3_214)
         );
  DFF_X1 tempStoreData_reg_213_ ( .D(U57_Z_213), .CK(clock), .Q(U6_DATA3_213)
         );
  DFF_X1 tempStoreData_reg_212_ ( .D(U57_Z_212), .CK(clock), .Q(U6_DATA3_212)
         );
  DFF_X1 tempStoreData_reg_211_ ( .D(U57_Z_211), .CK(clock), .Q(U6_DATA3_211)
         );
  DFF_X1 tempStoreData_reg_210_ ( .D(U57_Z_210), .CK(clock), .Q(U6_DATA3_210)
         );
  DFF_X1 tempStoreData_reg_209_ ( .D(U57_Z_209), .CK(clock), .Q(U6_DATA3_209)
         );
  DFF_X1 tempStoreData_reg_208_ ( .D(U57_Z_208), .CK(clock), .Q(U6_DATA3_208)
         );
  DFF_X1 tempStoreData_reg_207_ ( .D(U57_Z_207), .CK(clock), .Q(U6_DATA3_207)
         );
  DFF_X1 tempStoreData_reg_206_ ( .D(U57_Z_206), .CK(clock), .Q(U6_DATA3_206)
         );
  DFF_X1 tempStoreData_reg_205_ ( .D(U57_Z_205), .CK(clock), .Q(U6_DATA3_205)
         );
  DFF_X1 tempStoreData_reg_204_ ( .D(U57_Z_204), .CK(clock), .Q(U6_DATA3_204)
         );
  DFF_X1 tempStoreData_reg_203_ ( .D(U57_Z_203), .CK(clock), .Q(U6_DATA3_203)
         );
  DFF_X1 tempStoreData_reg_202_ ( .D(U57_Z_202), .CK(clock), .Q(U6_DATA3_202)
         );
  DFF_X1 tempStoreData_reg_201_ ( .D(U57_Z_201), .CK(clock), .Q(U6_DATA3_201)
         );
  DFF_X1 tempStoreData_reg_200_ ( .D(U57_Z_200), .CK(clock), .Q(U6_DATA3_200)
         );
  DFF_X1 tempStoreData_reg_199_ ( .D(U57_Z_199), .CK(clock), .Q(U6_DATA3_199)
         );
  DFF_X1 tempStoreData_reg_198_ ( .D(U57_Z_198), .CK(clock), .Q(U6_DATA3_198)
         );
  DFF_X1 tempStoreData_reg_197_ ( .D(U57_Z_197), .CK(clock), .Q(U6_DATA3_197)
         );
  DFF_X1 tempStoreData_reg_196_ ( .D(U57_Z_196), .CK(clock), .Q(U6_DATA3_196)
         );
  DFF_X1 tempStoreData_reg_195_ ( .D(U57_Z_195), .CK(clock), .Q(U6_DATA3_195)
         );
  DFF_X1 tempStoreData_reg_194_ ( .D(U57_Z_194), .CK(clock), .Q(U6_DATA3_194)
         );
  DFF_X1 tempStoreData_reg_193_ ( .D(U57_Z_193), .CK(clock), .Q(U6_DATA3_193)
         );
  DFF_X1 tempStoreData_reg_192_ ( .D(U57_Z_192), .CK(clock), .Q(U6_DATA3_192)
         );
  DFF_X2 tempStoreData_reg_175_ ( .D(U57_Z_175), .CK(clock), .QN(n126) );
  DFF_X2 tempStoreData_reg_174_ ( .D(U57_Z_174), .CK(clock), .QN(n127) );
  DFF_X2 tempStoreData_reg_173_ ( .D(U57_Z_173), .CK(clock), .QN(n128) );
  DFF_X2 tempStoreData_reg_172_ ( .D(U57_Z_172), .CK(clock), .QN(n129) );
  DFF_X2 tempStoreData_reg_171_ ( .D(U57_Z_171), .CK(clock), .QN(n130) );
  DFF_X2 tempStoreData_reg_170_ ( .D(U57_Z_170), .CK(clock), .QN(n131) );
  DFF_X2 tempStoreData_reg_169_ ( .D(U57_Z_169), .CK(clock), .QN(n132) );
  DFF_X2 tempStoreData_reg_168_ ( .D(U57_Z_168), .CK(clock), .QN(n133) );
  DFF_X2 tempStoreData_reg_167_ ( .D(U57_Z_167), .CK(clock), .QN(n134) );
  DFF_X2 tempStoreData_reg_166_ ( .D(U57_Z_166), .CK(clock), .QN(n135) );
  DFF_X2 tempStoreData_reg_165_ ( .D(U57_Z_165), .CK(clock), .QN(n136) );
  DFF_X2 tempStoreData_reg_164_ ( .D(U57_Z_164), .CK(clock), .QN(n137) );
  DFF_X2 tempStoreData_reg_163_ ( .D(U57_Z_163), .CK(clock), .QN(n138) );
  DFF_X2 tempStoreData_reg_162_ ( .D(U57_Z_162), .CK(clock), .QN(n139) );
  DFF_X2 tempStoreData_reg_161_ ( .D(U57_Z_161), .CK(clock), .QN(n140) );
  DFF_X2 tempStoreData_reg_160_ ( .D(U57_Z_160), .CK(clock), .QN(n141) );
  DFF_X2 tempStoreData_reg_159_ ( .D(U57_Z_159), .CK(clock), .QN(n142) );
  DFF_X2 tempStoreData_reg_158_ ( .D(U57_Z_158), .CK(clock), .QN(n143) );
  DFF_X2 tempStoreData_reg_157_ ( .D(U57_Z_157), .CK(clock), .QN(n144) );
  DFF_X2 tempStoreData_reg_156_ ( .D(U57_Z_156), .CK(clock), .QN(n145) );
  DFF_X2 tempStoreData_reg_155_ ( .D(U57_Z_155), .CK(clock), .QN(n146) );
  DFF_X2 tempStoreData_reg_154_ ( .D(U57_Z_154), .CK(clock), .QN(n147) );
  DFF_X2 tempStoreData_reg_153_ ( .D(U57_Z_153), .CK(clock), .QN(n148) );
  DFF_X2 tempStoreData_reg_152_ ( .D(U57_Z_152), .CK(clock), .QN(n149) );
  DFF_X2 tempStoreData_reg_151_ ( .D(U57_Z_151), .CK(clock), .QN(n150) );
  DFF_X2 tempStoreData_reg_150_ ( .D(U57_Z_150), .CK(clock), .QN(n151) );
  DFF_X2 tempStoreData_reg_149_ ( .D(U57_Z_149), .CK(clock), .QN(n152) );
  DFF_X2 tempStoreData_reg_148_ ( .D(U57_Z_148), .CK(clock), .QN(n153) );
  DFF_X2 tempStoreData_reg_147_ ( .D(U57_Z_147), .CK(clock), .QN(n154) );
  DFF_X2 tempStoreData_reg_146_ ( .D(U57_Z_146), .CK(clock), .QN(n155) );
  DFF_X2 tempStoreData_reg_145_ ( .D(U57_Z_145), .CK(clock), .QN(n156) );
  DFF_X2 tempStoreData_reg_144_ ( .D(U57_Z_144), .CK(clock), .QN(n157) );
  DFF_X2 tempStoreData_reg_143_ ( .D(U57_Z_143), .CK(clock), .QN(n158) );
  DFF_X2 tempStoreData_reg_142_ ( .D(U57_Z_142), .CK(clock), .QN(n159) );
  DFF_X2 tempStoreData_reg_141_ ( .D(U57_Z_141), .CK(clock), .QN(n160) );
  DFF_X2 tempStoreData_reg_140_ ( .D(U57_Z_140), .CK(clock), .QN(n161) );
  DFF_X2 tempStoreData_reg_139_ ( .D(U57_Z_139), .CK(clock), .QN(n162) );
  DFF_X2 tempStoreData_reg_138_ ( .D(U57_Z_138), .CK(clock), .QN(n163) );
  DFF_X2 tempStoreData_reg_137_ ( .D(U57_Z_137), .CK(clock), .QN(n164) );
  DFF_X2 tempStoreData_reg_136_ ( .D(U57_Z_136), .CK(clock), .QN(n165) );
  DFF_X2 tempStoreData_reg_135_ ( .D(U57_Z_135), .CK(clock), .QN(n166) );
  DFF_X2 tempStoreData_reg_134_ ( .D(U57_Z_134), .CK(clock), .QN(n167) );
  DFF_X2 tempStoreData_reg_133_ ( .D(U57_Z_133), .CK(clock), .QN(n168) );
  DFF_X2 tempStoreData_reg_132_ ( .D(U57_Z_132), .CK(clock), .QN(n169) );
  DFF_X2 tempStoreData_reg_131_ ( .D(U57_Z_131), .CK(clock), .QN(n170) );
  DFF_X2 tempStoreData_reg_130_ ( .D(U57_Z_130), .CK(clock), .QN(n171) );
  DFF_X2 tempStoreData_reg_129_ ( .D(U57_Z_129), .CK(clock), .QN(n172) );
  DFF_X2 tempStoreData_reg_128_ ( .D(U57_Z_128), .CK(clock), .QN(n173) );
  DFF_X2 tempStoreData_reg_99_ ( .D(U57_Z_99), .CK(clock), .QN(n186) );
  DFF_X2 tempStoreData_reg_98_ ( .D(U57_Z_98), .CK(clock), .QN(n187) );
  DFF_X2 tempStoreData_reg_97_ ( .D(U57_Z_97), .CK(clock), .QN(n188) );
  DFF_X2 tempStoreData_reg_96_ ( .D(U57_Z_96), .CK(clock), .QN(n189) );
  DFF_X2 tempStoreData_reg_95_ ( .D(U57_Z_95), .CK(clock), .QN(n190) );
  DFF_X2 tempStoreData_reg_94_ ( .D(U57_Z_94), .CK(clock), .QN(n191) );
  DFF_X2 tempStoreData_reg_93_ ( .D(U57_Z_93), .CK(clock), .QN(n192) );
  DFF_X2 tempStoreData_reg_92_ ( .D(U57_Z_92), .CK(clock), .QN(n193) );
  DFF_X2 tempStoreData_reg_91_ ( .D(U57_Z_91), .CK(clock), .QN(n194) );
  DFF_X2 tempStoreData_reg_90_ ( .D(U57_Z_90), .CK(clock), .QN(n195) );
  DFF_X2 tempStoreData_reg_89_ ( .D(U57_Z_89), .CK(clock), .QN(n196) );
  DFF_X2 tempStoreData_reg_88_ ( .D(U57_Z_88), .CK(clock), .QN(n197) );
  DFF_X2 tempStoreData_reg_87_ ( .D(U57_Z_87), .CK(clock), .QN(n198) );
  DFF_X2 tempStoreData_reg_86_ ( .D(U57_Z_86), .CK(clock), .QN(n199) );
  DFF_X2 tempStoreData_reg_85_ ( .D(U57_Z_85), .CK(clock), .QN(n200) );
  DFF_X2 tempStoreData_reg_84_ ( .D(U57_Z_84), .CK(clock), .QN(n201) );
  DFF_X2 tempStoreData_reg_83_ ( .D(U57_Z_83), .CK(clock), .QN(n202) );
  DFF_X2 tempStoreData_reg_82_ ( .D(U57_Z_82), .CK(clock), .QN(n203) );
  DFF_X2 tempStoreData_reg_81_ ( .D(U57_Z_81), .CK(clock), .QN(n204) );
  DFF_X2 tempStoreData_reg_80_ ( .D(U57_Z_80), .CK(clock), .QN(n205) );
  DFF_X2 tempStoreData_reg_79_ ( .D(U57_Z_79), .CK(clock), .QN(n206) );
  DFF_X2 tempStoreData_reg_78_ ( .D(U57_Z_78), .CK(clock), .QN(n207) );
  DFF_X2 tempStoreData_reg_77_ ( .D(U57_Z_77), .CK(clock), .QN(n208) );
  DFF_X2 tempStoreData_reg_76_ ( .D(U57_Z_76), .CK(clock), .QN(n209) );
  DFF_X2 tempStoreData_reg_75_ ( .D(U57_Z_75), .CK(clock), .QN(n210) );
  DFF_X2 tempStoreData_reg_74_ ( .D(U57_Z_74), .CK(clock), .QN(n211) );
  DFF_X2 tempStoreData_reg_73_ ( .D(U57_Z_73), .CK(clock), .QN(n212) );
  DFF_X2 tempStoreData_reg_72_ ( .D(U57_Z_72), .CK(clock), .QN(n213) );
  DFF_X2 tempStoreData_reg_71_ ( .D(U57_Z_71), .CK(clock), .QN(n214) );
  DFF_X2 tempStoreData_reg_70_ ( .D(U57_Z_70), .CK(clock), .QN(n215) );
  DFF_X2 tempStoreData_reg_69_ ( .D(U57_Z_69), .CK(clock), .QN(n216) );
  DFF_X2 tempStoreData_reg_68_ ( .D(U57_Z_68), .CK(clock), .QN(n217) );
  DFF_X2 tempStoreData_reg_67_ ( .D(U57_Z_67), .CK(clock), .QN(n218) );
  DFF_X2 tempStoreData_reg_66_ ( .D(U57_Z_66), .CK(clock), .QN(n219) );
  DFF_X2 tempStoreData_reg_65_ ( .D(U57_Z_65), .CK(clock), .QN(n220) );
  DFF_X2 tempStoreData_reg_64_ ( .D(U57_Z_64), .CK(clock), .QN(n221) );
  DFF_X2 tempStoreData_reg_111_ ( .D(U57_Z_111), .CK(clock), .QN(n174) );
  DFF_X2 tempStoreData_reg_110_ ( .D(U57_Z_110), .CK(clock), .QN(n175) );
  DFF_X2 tempStoreData_reg_109_ ( .D(U57_Z_109), .CK(clock), .QN(n176) );
  DFF_X2 tempStoreData_reg_108_ ( .D(U57_Z_108), .CK(clock), .QN(n177) );
  DFF_X2 tempStoreData_reg_107_ ( .D(U57_Z_107), .CK(clock), .QN(n178) );
  DFF_X2 tempStoreData_reg_106_ ( .D(U57_Z_106), .CK(clock), .QN(n179) );
  DFF_X2 tempStoreData_reg_105_ ( .D(U57_Z_105), .CK(clock), .QN(n180) );
  DFF_X2 tempStoreData_reg_104_ ( .D(U57_Z_104), .CK(clock), .QN(n181) );
  DFF_X2 tempStoreData_reg_103_ ( .D(U57_Z_103), .CK(clock), .QN(n182) );
  DFF_X2 tempStoreData_reg_102_ ( .D(U57_Z_102), .CK(clock), .QN(n183) );
  DFF_X2 tempStoreData_reg_101_ ( .D(U57_Z_101), .CK(clock), .QN(n184) );
  DFF_X2 tempStoreData_reg_100_ ( .D(U57_Z_100), .CK(clock), .QN(n185) );
  DFF_X1 tempStoreData_reg_63_ ( .D(U57_Z_63), .CK(clock), .Q(U6_DATA3_63) );
  DFF_X1 op_writeData_reg_63_ ( .D(n118), .CK(clock), .Q(op_writeData[63]) );
  DFF_X1 tempStoreData_reg_62_ ( .D(U57_Z_62), .CK(clock), .Q(U6_DATA3_62) );
  DFF_X1 op_writeData_reg_62_ ( .D(n117), .CK(clock), .Q(op_writeData[62]) );
  DFF_X1 tempStoreData_reg_61_ ( .D(U57_Z_61), .CK(clock), .Q(U6_DATA3_61) );
  DFF_X1 op_writeData_reg_61_ ( .D(n116), .CK(clock), .Q(op_writeData[61]) );
  DFF_X1 tempStoreData_reg_60_ ( .D(U57_Z_60), .CK(clock), .Q(U6_DATA3_60) );
  DFF_X1 op_writeData_reg_60_ ( .D(n115), .CK(clock), .Q(op_writeData[60]) );
  DFF_X1 tempStoreData_reg_59_ ( .D(U57_Z_59), .CK(clock), .Q(U6_DATA3_59) );
  DFF_X1 op_writeData_reg_59_ ( .D(n114), .CK(clock), .Q(op_writeData[59]) );
  DFF_X1 tempStoreData_reg_58_ ( .D(U57_Z_58), .CK(clock), .Q(U6_DATA3_58) );
  DFF_X1 op_writeData_reg_58_ ( .D(n113), .CK(clock), .Q(op_writeData[58]) );
  DFF_X1 tempStoreData_reg_57_ ( .D(U57_Z_57), .CK(clock), .Q(U6_DATA3_57) );
  DFF_X1 op_writeData_reg_57_ ( .D(n112), .CK(clock), .Q(op_writeData[57]) );
  DFF_X1 tempStoreData_reg_56_ ( .D(U57_Z_56), .CK(clock), .Q(U6_DATA3_56) );
  DFF_X1 op_writeData_reg_56_ ( .D(n111), .CK(clock), .Q(op_writeData[56]) );
  DFF_X1 tempStoreData_reg_55_ ( .D(U57_Z_55), .CK(clock), .Q(U6_DATA3_55) );
  DFF_X1 op_writeData_reg_55_ ( .D(n110), .CK(clock), .Q(op_writeData[55]) );
  DFF_X1 tempStoreData_reg_54_ ( .D(U57_Z_54), .CK(clock), .Q(U6_DATA3_54) );
  DFF_X1 op_writeData_reg_54_ ( .D(n109), .CK(clock), .Q(op_writeData[54]) );
  DFF_X1 tempStoreData_reg_53_ ( .D(U57_Z_53), .CK(clock), .Q(U6_DATA3_53) );
  DFF_X1 op_writeData_reg_53_ ( .D(n108), .CK(clock), .Q(op_writeData[53]) );
  DFF_X1 tempStoreData_reg_52_ ( .D(U57_Z_52), .CK(clock), .Q(U6_DATA3_52) );
  DFF_X1 op_writeData_reg_52_ ( .D(n107), .CK(clock), .Q(op_writeData[52]) );
  DFF_X1 tempStoreData_reg_51_ ( .D(U57_Z_51), .CK(clock), .Q(U6_DATA3_51) );
  DFF_X1 op_writeData_reg_51_ ( .D(n106), .CK(clock), .Q(op_writeData[51]) );
  DFF_X1 tempStoreData_reg_50_ ( .D(U57_Z_50), .CK(clock), .Q(U6_DATA3_50) );
  DFF_X1 op_writeData_reg_50_ ( .D(n105), .CK(clock), .Q(op_writeData[50]) );
  DFF_X1 tempStoreData_reg_49_ ( .D(U57_Z_49), .CK(clock), .Q(U6_DATA3_49) );
  DFF_X1 op_writeData_reg_49_ ( .D(n104), .CK(clock), .Q(op_writeData[49]) );
  DFF_X1 tempStoreData_reg_48_ ( .D(U57_Z_48), .CK(clock), .Q(U6_DATA3_48) );
  DFF_X1 op_writeData_reg_48_ ( .D(n103), .CK(clock), .Q(op_writeData[48]) );
  DFF_X1 tempStoreData_reg_255_ ( .D(U57_Z_255), .CK(clock), .Q(U6_DATA3_255)
         );
  DFF_X1 op_writeData_reg_255_ ( .D(n102), .CK(clock), .Q(op_writeData[255])
         );
  DFF_X1 tempStoreData_reg_254_ ( .D(U57_Z_254), .CK(clock), .Q(U6_DATA3_254)
         );
  DFF_X1 op_writeData_reg_254_ ( .D(n101), .CK(clock), .Q(op_writeData[254])
         );
  DFF_X1 tempStoreData_reg_253_ ( .D(U57_Z_253), .CK(clock), .Q(U6_DATA3_253)
         );
  DFF_X1 op_writeData_reg_253_ ( .D(n100), .CK(clock), .Q(op_writeData[253])
         );
  DFF_X1 tempStoreData_reg_252_ ( .D(U57_Z_252), .CK(clock), .Q(U6_DATA3_252)
         );
  DFF_X1 op_writeData_reg_252_ ( .D(n99), .CK(clock), .Q(op_writeData[252]) );
  DFF_X1 tempStoreData_reg_251_ ( .D(U57_Z_251), .CK(clock), .Q(U6_DATA3_251)
         );
  DFF_X1 op_writeData_reg_251_ ( .D(n98), .CK(clock), .Q(op_writeData[251]) );
  DFF_X1 tempStoreData_reg_250_ ( .D(U57_Z_250), .CK(clock), .Q(U6_DATA3_250)
         );
  DFF_X1 op_writeData_reg_250_ ( .D(n97), .CK(clock), .Q(op_writeData[250]) );
  DFF_X1 tempStoreData_reg_249_ ( .D(U57_Z_249), .CK(clock), .Q(U6_DATA3_249)
         );
  DFF_X1 op_writeData_reg_249_ ( .D(n96), .CK(clock), .Q(op_writeData[249]) );
  DFF_X1 tempStoreData_reg_248_ ( .D(U57_Z_248), .CK(clock), .Q(U6_DATA3_248)
         );
  DFF_X1 op_writeData_reg_248_ ( .D(n95), .CK(clock), .Q(op_writeData[248]) );
  DFF_X1 tempStoreData_reg_247_ ( .D(U57_Z_247), .CK(clock), .Q(U6_DATA3_247)
         );
  DFF_X1 op_writeData_reg_247_ ( .D(n94), .CK(clock), .Q(op_writeData[247]) );
  DFF_X1 tempStoreData_reg_246_ ( .D(U57_Z_246), .CK(clock), .Q(U6_DATA3_246)
         );
  DFF_X1 op_writeData_reg_246_ ( .D(n93), .CK(clock), .Q(op_writeData[246]) );
  DFF_X1 tempStoreData_reg_245_ ( .D(U57_Z_245), .CK(clock), .Q(U6_DATA3_245)
         );
  DFF_X1 op_writeData_reg_245_ ( .D(n92), .CK(clock), .Q(op_writeData[245]) );
  DFF_X1 tempStoreData_reg_244_ ( .D(U57_Z_244), .CK(clock), .Q(U6_DATA3_244)
         );
  DFF_X1 op_writeData_reg_244_ ( .D(n91), .CK(clock), .Q(op_writeData[244]) );
  DFF_X1 tempStoreData_reg_243_ ( .D(U57_Z_243), .CK(clock), .Q(U6_DATA3_243)
         );
  DFF_X1 op_writeData_reg_243_ ( .D(n90), .CK(clock), .Q(op_writeData[243]) );
  DFF_X1 tempStoreData_reg_242_ ( .D(U57_Z_242), .CK(clock), .Q(U6_DATA3_242)
         );
  DFF_X1 op_writeData_reg_242_ ( .D(n89), .CK(clock), .Q(op_writeData[242]) );
  DFF_X1 tempStoreData_reg_241_ ( .D(U57_Z_241), .CK(clock), .Q(U6_DATA3_241)
         );
  DFF_X1 op_writeData_reg_241_ ( .D(n88), .CK(clock), .Q(op_writeData[241]) );
  DFF_X1 tempStoreData_reg_240_ ( .D(U57_Z_240), .CK(clock), .Q(U6_DATA3_240)
         );
  DFF_X1 op_writeData_reg_240_ ( .D(n87), .CK(clock), .Q(op_writeData[240]) );
  DFF_X1 tempStoreData_reg_191_ ( .D(U57_Z_191), .CK(clock), .Q(U6_DATA3_191)
         );
  DFF_X1 op_writeData_reg_191_ ( .D(n38), .CK(clock), .Q(op_writeData[191]) );
  DFF_X1 tempStoreData_reg_190_ ( .D(U57_Z_190), .CK(clock), .Q(U6_DATA3_190)
         );
  DFF_X1 op_writeData_reg_190_ ( .D(n37), .CK(clock), .Q(op_writeData[190]) );
  DFF_X1 tempStoreData_reg_189_ ( .D(U57_Z_189), .CK(clock), .Q(U6_DATA3_189)
         );
  DFF_X1 op_writeData_reg_189_ ( .D(n36), .CK(clock), .Q(op_writeData[189]) );
  DFF_X1 tempStoreData_reg_188_ ( .D(U57_Z_188), .CK(clock), .Q(U6_DATA3_188)
         );
  DFF_X1 op_writeData_reg_188_ ( .D(n35), .CK(clock), .Q(op_writeData[188]) );
  DFF_X1 tempStoreData_reg_187_ ( .D(U57_Z_187), .CK(clock), .Q(U6_DATA3_187)
         );
  DFF_X1 op_writeData_reg_187_ ( .D(n34), .CK(clock), .Q(op_writeData[187]) );
  DFF_X1 tempStoreData_reg_186_ ( .D(U57_Z_186), .CK(clock), .Q(U6_DATA3_186)
         );
  DFF_X1 op_writeData_reg_186_ ( .D(n33), .CK(clock), .Q(op_writeData[186]) );
  DFF_X1 tempStoreData_reg_185_ ( .D(U57_Z_185), .CK(clock), .Q(U6_DATA3_185)
         );
  DFF_X1 op_writeData_reg_185_ ( .D(n32), .CK(clock), .Q(op_writeData[185]) );
  DFF_X1 tempStoreData_reg_184_ ( .D(U57_Z_184), .CK(clock), .Q(U6_DATA3_184)
         );
  DFF_X1 op_writeData_reg_184_ ( .D(n31), .CK(clock), .Q(op_writeData[184]) );
  DFF_X1 tempStoreData_reg_183_ ( .D(U57_Z_183), .CK(clock), .Q(U6_DATA3_183)
         );
  DFF_X1 op_writeData_reg_183_ ( .D(n30), .CK(clock), .Q(op_writeData[183]) );
  DFF_X1 tempStoreData_reg_182_ ( .D(U57_Z_182), .CK(clock), .Q(U6_DATA3_182)
         );
  DFF_X1 op_writeData_reg_182_ ( .D(n29), .CK(clock), .Q(op_writeData[182]) );
  DFF_X1 tempStoreData_reg_181_ ( .D(U57_Z_181), .CK(clock), .Q(U6_DATA3_181)
         );
  DFF_X1 op_writeData_reg_181_ ( .D(n28), .CK(clock), .Q(op_writeData[181]) );
  DFF_X1 tempStoreData_reg_180_ ( .D(U57_Z_180), .CK(clock), .Q(U6_DATA3_180)
         );
  DFF_X1 op_writeData_reg_180_ ( .D(n27), .CK(clock), .Q(op_writeData[180]) );
  DFF_X1 tempStoreData_reg_179_ ( .D(U57_Z_179), .CK(clock), .Q(U6_DATA3_179)
         );
  DFF_X1 op_writeData_reg_179_ ( .D(n26), .CK(clock), .Q(op_writeData[179]) );
  DFF_X1 tempStoreData_reg_178_ ( .D(U57_Z_178), .CK(clock), .Q(U6_DATA3_178)
         );
  DFF_X1 op_writeData_reg_178_ ( .D(n25), .CK(clock), .Q(op_writeData[178]) );
  DFF_X1 tempStoreData_reg_177_ ( .D(U57_Z_177), .CK(clock), .Q(U6_DATA3_177)
         );
  DFF_X1 op_writeData_reg_177_ ( .D(n24), .CK(clock), .Q(op_writeData[177]) );
  DFF_X1 tempStoreData_reg_176_ ( .D(U57_Z_176), .CK(clock), .Q(U6_DATA3_176)
         );
  DFF_X1 op_writeData_reg_176_ ( .D(n23), .CK(clock), .Q(op_writeData[176]) );
  DFF_X1 tempStoreData_reg_127_ ( .D(U57_Z_127), .CK(clock), .Q(U6_DATA3_127)
         );
  DFF_X1 op_writeData_reg_127_ ( .D(n22), .CK(clock), .Q(op_writeData[127]) );
  DFF_X1 tempStoreData_reg_126_ ( .D(U57_Z_126), .CK(clock), .Q(U6_DATA3_126)
         );
  DFF_X1 op_writeData_reg_126_ ( .D(n21), .CK(clock), .Q(op_writeData[126]) );
  DFF_X1 tempStoreData_reg_125_ ( .D(U57_Z_125), .CK(clock), .Q(U6_DATA3_125)
         );
  DFF_X1 op_writeData_reg_125_ ( .D(n20), .CK(clock), .Q(op_writeData[125]) );
  DFF_X1 tempStoreData_reg_124_ ( .D(U57_Z_124), .CK(clock), .Q(U6_DATA3_124)
         );
  DFF_X1 op_writeData_reg_124_ ( .D(n19), .CK(clock), .Q(op_writeData[124]) );
  DFF_X1 tempStoreData_reg_123_ ( .D(U57_Z_123), .CK(clock), .Q(U6_DATA3_123)
         );
  DFF_X1 op_writeData_reg_123_ ( .D(n18), .CK(clock), .Q(op_writeData[123]) );
  DFF_X1 tempStoreData_reg_122_ ( .D(U57_Z_122), .CK(clock), .Q(U6_DATA3_122)
         );
  DFF_X1 op_writeData_reg_122_ ( .D(n17), .CK(clock), .Q(op_writeData[122]) );
  DFF_X1 tempStoreData_reg_121_ ( .D(U57_Z_121), .CK(clock), .Q(U6_DATA3_121)
         );
  DFF_X1 op_writeData_reg_121_ ( .D(n16), .CK(clock), .Q(op_writeData[121]) );
  DFF_X1 tempStoreData_reg_120_ ( .D(U57_Z_120), .CK(clock), .Q(U6_DATA3_120)
         );
  DFF_X1 op_writeData_reg_120_ ( .D(n15), .CK(clock), .Q(op_writeData[120]) );
  DFF_X1 tempStoreData_reg_119_ ( .D(U57_Z_119), .CK(clock), .Q(U6_DATA3_119)
         );
  DFF_X1 op_writeData_reg_119_ ( .D(n14), .CK(clock), .Q(op_writeData[119]) );
  DFF_X1 tempStoreData_reg_118_ ( .D(U57_Z_118), .CK(clock), .Q(U6_DATA3_118)
         );
  DFF_X1 op_writeData_reg_118_ ( .D(n13), .CK(clock), .Q(op_writeData[118]) );
  DFF_X1 tempStoreData_reg_117_ ( .D(U57_Z_117), .CK(clock), .Q(U6_DATA3_117)
         );
  DFF_X1 op_writeData_reg_117_ ( .D(n12), .CK(clock), .Q(op_writeData[117]) );
  DFF_X1 tempStoreData_reg_116_ ( .D(U57_Z_116), .CK(clock), .Q(U6_DATA3_116)
         );
  DFF_X1 op_writeData_reg_116_ ( .D(n11), .CK(clock), .Q(op_writeData[116]) );
  DFF_X1 tempStoreData_reg_115_ ( .D(U57_Z_115), .CK(clock), .Q(U6_DATA3_115)
         );
  DFF_X1 op_writeData_reg_115_ ( .D(n10), .CK(clock), .Q(op_writeData[115]) );
  DFF_X1 tempStoreData_reg_114_ ( .D(U57_Z_114), .CK(clock), .Q(U6_DATA3_114)
         );
  DFF_X1 op_writeData_reg_114_ ( .D(n9), .CK(clock), .Q(op_writeData[114]) );
  DFF_X1 tempStoreData_reg_113_ ( .D(U57_Z_113), .CK(clock), .Q(U6_DATA3_113)
         );
  DFF_X1 op_writeData_reg_113_ ( .D(n8), .CK(clock), .Q(op_writeData[113]) );
  DFF_X1 tempStoreData_reg_112_ ( .D(U57_Z_112), .CK(clock), .Q(U6_DATA3_112)
         );
  DFF_X1 op_writeData_reg_112_ ( .D(n7), .CK(clock), .Q(op_writeData[112]) );
  DFF_X2 tempStoreData_reg_9_ ( .D(U57_Z_9), .CK(clock), .QN(n260) );
  DFF_X2 tempStoreData_reg_8_ ( .D(U57_Z_8), .CK(clock), .QN(n261) );
  DFF_X2 tempStoreData_reg_7_ ( .D(U57_Z_7), .CK(clock), .QN(n262) );
  DFF_X2 tempStoreData_reg_6_ ( .D(U57_Z_6), .CK(clock), .QN(n263) );
  DFF_X2 tempStoreData_reg_5_ ( .D(U57_Z_5), .CK(clock), .QN(n264) );
  DFF_X2 tempStoreData_reg_47_ ( .D(U57_Z_47), .CK(clock), .QN(n222) );
  DFF_X2 tempStoreData_reg_46_ ( .D(U57_Z_46), .CK(clock), .QN(n223) );
  DFF_X2 tempStoreData_reg_45_ ( .D(U57_Z_45), .CK(clock), .QN(n224) );
  DFF_X2 tempStoreData_reg_44_ ( .D(U57_Z_44), .CK(clock), .QN(n225) );
  DFF_X2 tempStoreData_reg_43_ ( .D(U57_Z_43), .CK(clock), .QN(n226) );
  DFF_X2 tempStoreData_reg_42_ ( .D(U57_Z_42), .CK(clock), .QN(n227) );
  DFF_X2 tempStoreData_reg_41_ ( .D(U57_Z_41), .CK(clock), .QN(n228) );
  DFF_X2 tempStoreData_reg_40_ ( .D(U57_Z_40), .CK(clock), .QN(n229) );
  DFF_X2 tempStoreData_reg_4_ ( .D(U57_Z_4), .CK(clock), .QN(n265) );
  DFF_X2 tempStoreData_reg_39_ ( .D(U57_Z_39), .CK(clock), .QN(n230) );
  DFF_X2 tempStoreData_reg_38_ ( .D(U57_Z_38), .CK(clock), .QN(n231) );
  DFF_X2 tempStoreData_reg_37_ ( .D(U57_Z_37), .CK(clock), .QN(n232) );
  DFF_X2 tempStoreData_reg_36_ ( .D(U57_Z_36), .CK(clock), .QN(n233) );
  DFF_X2 tempStoreData_reg_35_ ( .D(U57_Z_35), .CK(clock), .QN(n234) );
  DFF_X2 tempStoreData_reg_34_ ( .D(U57_Z_34), .CK(clock), .QN(n235) );
  DFF_X2 tempStoreData_reg_33_ ( .D(U57_Z_33), .CK(clock), .QN(n236) );
  DFF_X2 tempStoreData_reg_32_ ( .D(U57_Z_32), .CK(clock), .QN(n237) );
  DFF_X2 tempStoreData_reg_31_ ( .D(U57_Z_31), .CK(clock), .QN(n238) );
  DFF_X2 tempStoreData_reg_30_ ( .D(U57_Z_30), .CK(clock), .QN(n239) );
  DFF_X2 tempStoreData_reg_3_ ( .D(U57_Z_3), .CK(clock), .QN(n266) );
  DFF_X2 tempStoreData_reg_29_ ( .D(U57_Z_29), .CK(clock), .QN(n240) );
  DFF_X2 tempStoreData_reg_28_ ( .D(U57_Z_28), .CK(clock), .QN(n241) );
  DFF_X2 tempStoreData_reg_27_ ( .D(U57_Z_27), .CK(clock), .QN(n242) );
  DFF_X2 tempStoreData_reg_26_ ( .D(U57_Z_26), .CK(clock), .QN(n243) );
  DFF_X2 tempStoreData_reg_25_ ( .D(U57_Z_25), .CK(clock), .QN(n244) );
  DFF_X2 tempStoreData_reg_24_ ( .D(U57_Z_24), .CK(clock), .QN(n245) );
  DFF_X2 tempStoreData_reg_23_ ( .D(U57_Z_23), .CK(clock), .QN(n246) );
  DFF_X2 tempStoreData_reg_22_ ( .D(U57_Z_22), .CK(clock), .QN(n247) );
  DFF_X2 tempStoreData_reg_21_ ( .D(U57_Z_21), .CK(clock), .QN(n248) );
  DFF_X2 tempStoreData_reg_20_ ( .D(U57_Z_20), .CK(clock), .QN(n249) );
  DFF_X2 tempStoreData_reg_2_ ( .D(U57_Z_2), .CK(clock), .QN(n267) );
  DFF_X2 tempStoreData_reg_19_ ( .D(U57_Z_19), .CK(clock), .QN(n250) );
  DFF_X2 tempStoreData_reg_18_ ( .D(U57_Z_18), .CK(clock), .QN(n251) );
  DFF_X2 tempStoreData_reg_17_ ( .D(U57_Z_17), .CK(clock), .QN(n252) );
  DFF_X2 tempStoreData_reg_16_ ( .D(U57_Z_16), .CK(clock), .QN(n253) );
  DFF_X2 tempStoreData_reg_15_ ( .D(U57_Z_15), .CK(clock), .QN(n254) );
  DFF_X2 tempStoreData_reg_14_ ( .D(U57_Z_14), .CK(clock), .QN(n255) );
  DFF_X2 tempStoreData_reg_13_ ( .D(U57_Z_13), .CK(clock), .QN(n256) );
  DFF_X2 tempStoreData_reg_12_ ( .D(U57_Z_12), .CK(clock), .QN(n257) );
  DFF_X2 tempStoreData_reg_11_ ( .D(U57_Z_11), .CK(clock), .QN(n258) );
  DFF_X2 tempStoreData_reg_10_ ( .D(U57_Z_10), .CK(clock), .QN(n259) );
  DFF_X2 tempStoreData_reg_1_ ( .D(U57_Z_1), .CK(clock), .QN(n268) );
  DFF_X2 tempStoreData_reg_0_ ( .D(U57_Z_0), .CK(clock), .QN(n269) );
  DFF_X2 tempComputedDiagVal1_reg_47_ ( .D(n1323), .CK(clock), .QN(n347) );
  DFF_X2 tempComputedDiagVal1_reg_46_ ( .D(n1322), .CK(clock), .QN(n348) );
  DFF_X2 tempComputedDiagVal1_reg_45_ ( .D(n1321), .CK(clock), .QN(n349) );
  DFF_X2 tempComputedDiagVal1_reg_44_ ( .D(n1320), .CK(clock), .QN(n350) );
  DFF_X2 tempComputedDiagVal1_reg_43_ ( .D(n1319), .CK(clock), .QN(n351) );
  DFF_X2 tempComputedDiagVal1_reg_42_ ( .D(n1318), .CK(clock), .QN(n352) );
  DFF_X2 tempComputedDiagVal1_reg_41_ ( .D(n1317), .CK(clock), .QN(n353) );
  DFF_X2 tempComputedDiagVal1_reg_40_ ( .D(n1316), .CK(clock), .QN(n354) );
  DFF_X2 tempComputedDiagVal1_reg_39_ ( .D(n1315), .CK(clock), .QN(n355) );
  DFF_X2 tempComputedDiagVal1_reg_38_ ( .D(n1314), .CK(clock), .QN(n356) );
  DFF_X2 tempComputedDiagVal1_reg_37_ ( .D(n1313), .CK(clock), .QN(n357) );
  DFF_X2 tempComputedDiagVal1_reg_36_ ( .D(n1312), .CK(clock), .QN(n358) );
  DFF_X2 tempComputedDiagVal1_reg_35_ ( .D(n1311), .CK(clock), .QN(n359) );
  DFF_X2 tempComputedDiagVal1_reg_34_ ( .D(n1310), .CK(clock), .QN(n360) );
  DFF_X2 tempComputedDiagVal1_reg_33_ ( .D(n1309), .CK(clock), .QN(n361) );
  DFF_X2 tempComputedDiagVal1_reg_32_ ( .D(n1308), .CK(clock), .QN(n362) );
  DFF_X2 tempComputedDiagVal1_reg_31_ ( .D(n1307), .CK(clock), .QN(n363) );
  DFF_X2 tempComputedDiagVal1_reg_30_ ( .D(n1306), .CK(clock), .QN(n364) );
  DFF_X2 tempComputedDiagVal1_reg_29_ ( .D(n1305), .CK(clock), .QN(n365) );
  DFF_X2 tempComputedDiagVal1_reg_28_ ( .D(n1304), .CK(clock), .QN(n366) );
  DFF_X2 tempComputedDiagVal1_reg_27_ ( .D(n1303), .CK(clock), .QN(n367) );
  DFF_X2 tempComputedDiagVal1_reg_26_ ( .D(n1302), .CK(clock), .QN(n368) );
  DFF_X2 tempComputedDiagVal1_reg_25_ ( .D(n1301), .CK(clock), .QN(n369) );
  DFF_X2 tempComputedDiagVal1_reg_24_ ( .D(n1300), .CK(clock), .QN(n370) );
  DFF_X2 tempComputedDiagVal1_reg_23_ ( .D(n1299), .CK(clock), .QN(n371) );
  DFF_X2 tempComputedDiagVal1_reg_22_ ( .D(n1298), .CK(clock), .QN(n372) );
  DFF_X2 tempComputedDiagVal1_reg_21_ ( .D(n1297), .CK(clock), .QN(n373) );
  DFF_X2 tempComputedDiagVal1_reg_20_ ( .D(n1296), .CK(clock), .QN(n374) );
  DFF_X2 tempComputedDiagVal1_reg_19_ ( .D(n1295), .CK(clock), .QN(n375) );
  DFF_X2 tempComputedDiagVal1_reg_18_ ( .D(n1294), .CK(clock), .QN(n376) );
  DFF_X2 tempComputedDiagVal1_reg_17_ ( .D(n1293), .CK(clock), .QN(n377) );
  DFF_X2 tempComputedDiagVal1_reg_16_ ( .D(n1292), .CK(clock), .QN(n378) );
  DFF_X2 tempComputedDiagVal1_reg_15_ ( .D(n1291), .CK(clock), .QN(n379) );
  DFF_X2 tempComputedDiagVal1_reg_14_ ( .D(n1290), .CK(clock), .QN(n380) );
  DFF_X2 tempComputedDiagVal1_reg_13_ ( .D(n1289), .CK(clock), .QN(n381) );
  DFF_X2 tempComputedDiagVal1_reg_12_ ( .D(n1288), .CK(clock), .QN(n382) );
  DFF_X2 tempComputedDiagVal1_reg_11_ ( .D(n1287), .CK(clock), .QN(n383) );
  DFF_X2 tempComputedDiagVal1_reg_10_ ( .D(n1286), .CK(clock), .QN(n384) );
  DFF_X2 tempComputedDiagVal1_reg_9_ ( .D(n1285), .CK(clock), .QN(n385) );
  DFF_X2 tempComputedDiagVal1_reg_8_ ( .D(n1284), .CK(clock), .QN(n386) );
  DFF_X2 tempComputedDiagVal1_reg_7_ ( .D(n1283), .CK(clock), .QN(n387) );
  DFF_X2 tempComputedDiagVal1_reg_6_ ( .D(n1282), .CK(clock), .QN(n388) );
  DFF_X2 tempComputedDiagVal1_reg_5_ ( .D(n1281), .CK(clock), .QN(n389) );
  DFF_X2 tempComputedDiagVal1_reg_4_ ( .D(n1280), .CK(clock), .QN(n390) );
  DFF_X2 tempComputedDiagVal1_reg_3_ ( .D(n1279), .CK(clock), .QN(n391) );
  DFF_X2 tempComputedDiagVal1_reg_2_ ( .D(n1278), .CK(clock), .QN(n392) );
  DFF_X2 tempComputedDiagVal1_reg_1_ ( .D(n1277), .CK(clock), .QN(n393) );
  DFF_X2 tempComputedDiagVal1_reg_0_ ( .D(n1276), .CK(clock), .QN(n394) );
  DFF_X2 tempComputedDiagVal2_reg_47_ ( .D(n1275), .CK(clock), .QN(n395) );
  DFF_X1 op_writeData_reg_47_ ( .D(U62_Z_47), .CK(clock), .Q(op_writeData[47])
         );
  DFF_X1 op_writeData_reg_239_ ( .D(n86), .CK(clock), .Q(op_writeData[239]) );
  DFF_X1 op_writeData_reg_175_ ( .D(U62_Z_175), .CK(clock), .Q(
        op_writeData[175]) );
  DFF_X1 op_writeData_reg_111_ ( .D(U62_Z_111), .CK(clock), .Q(
        op_writeData[111]) );
  DFF_X2 tempComputedDiagVal2_reg_46_ ( .D(n1274), .CK(clock), .QN(n396) );
  DFF_X1 op_writeData_reg_46_ ( .D(U62_Z_46), .CK(clock), .Q(op_writeData[46])
         );
  DFF_X1 op_writeData_reg_238_ ( .D(n85), .CK(clock), .Q(op_writeData[238]) );
  DFF_X1 op_writeData_reg_174_ ( .D(U62_Z_174), .CK(clock), .Q(
        op_writeData[174]) );
  DFF_X1 op_writeData_reg_110_ ( .D(U62_Z_110), .CK(clock), .Q(
        op_writeData[110]) );
  DFF_X2 tempComputedDiagVal2_reg_45_ ( .D(n1273), .CK(clock), .QN(n397) );
  DFF_X1 op_writeData_reg_45_ ( .D(U62_Z_45), .CK(clock), .Q(op_writeData[45])
         );
  DFF_X1 op_writeData_reg_237_ ( .D(n84), .CK(clock), .Q(op_writeData[237]) );
  DFF_X1 op_writeData_reg_173_ ( .D(U62_Z_173), .CK(clock), .Q(
        op_writeData[173]) );
  DFF_X1 op_writeData_reg_109_ ( .D(U62_Z_109), .CK(clock), .Q(
        op_writeData[109]) );
  DFF_X2 tempComputedDiagVal2_reg_44_ ( .D(n1272), .CK(clock), .QN(n398) );
  DFF_X1 op_writeData_reg_44_ ( .D(U62_Z_44), .CK(clock), .Q(op_writeData[44])
         );
  DFF_X1 op_writeData_reg_236_ ( .D(n83), .CK(clock), .Q(op_writeData[236]) );
  DFF_X1 op_writeData_reg_172_ ( .D(U62_Z_172), .CK(clock), .Q(
        op_writeData[172]) );
  DFF_X1 op_writeData_reg_108_ ( .D(U62_Z_108), .CK(clock), .Q(
        op_writeData[108]) );
  DFF_X2 tempComputedDiagVal2_reg_43_ ( .D(n1271), .CK(clock), .QN(n399) );
  DFF_X1 op_writeData_reg_43_ ( .D(U62_Z_43), .CK(clock), .Q(op_writeData[43])
         );
  DFF_X1 op_writeData_reg_235_ ( .D(n82), .CK(clock), .Q(op_writeData[235]) );
  DFF_X1 op_writeData_reg_171_ ( .D(U62_Z_171), .CK(clock), .Q(
        op_writeData[171]) );
  DFF_X1 op_writeData_reg_107_ ( .D(U62_Z_107), .CK(clock), .Q(
        op_writeData[107]) );
  DFF_X2 tempComputedDiagVal2_reg_42_ ( .D(n1270), .CK(clock), .QN(n400) );
  DFF_X1 op_writeData_reg_42_ ( .D(U62_Z_42), .CK(clock), .Q(op_writeData[42])
         );
  DFF_X1 op_writeData_reg_234_ ( .D(n81), .CK(clock), .Q(op_writeData[234]) );
  DFF_X1 op_writeData_reg_170_ ( .D(U62_Z_170), .CK(clock), .Q(
        op_writeData[170]) );
  DFF_X1 op_writeData_reg_106_ ( .D(U62_Z_106), .CK(clock), .Q(
        op_writeData[106]) );
  DFF_X2 tempComputedDiagVal2_reg_41_ ( .D(n1269), .CK(clock), .QN(n401) );
  DFF_X1 op_writeData_reg_41_ ( .D(U62_Z_41), .CK(clock), .Q(op_writeData[41])
         );
  DFF_X1 op_writeData_reg_233_ ( .D(n80), .CK(clock), .Q(op_writeData[233]) );
  DFF_X1 op_writeData_reg_169_ ( .D(U62_Z_169), .CK(clock), .Q(
        op_writeData[169]) );
  DFF_X1 op_writeData_reg_105_ ( .D(U62_Z_105), .CK(clock), .Q(
        op_writeData[105]) );
  DFF_X2 tempComputedDiagVal2_reg_40_ ( .D(n1268), .CK(clock), .QN(n402) );
  DFF_X1 op_writeData_reg_40_ ( .D(U62_Z_40), .CK(clock), .Q(op_writeData[40])
         );
  DFF_X1 op_writeData_reg_232_ ( .D(n79), .CK(clock), .Q(op_writeData[232]) );
  DFF_X1 op_writeData_reg_168_ ( .D(U62_Z_168), .CK(clock), .Q(
        op_writeData[168]) );
  DFF_X1 op_writeData_reg_104_ ( .D(U62_Z_104), .CK(clock), .Q(
        op_writeData[104]) );
  DFF_X2 tempComputedDiagVal2_reg_39_ ( .D(n1267), .CK(clock), .QN(n403) );
  DFF_X1 op_writeData_reg_39_ ( .D(U62_Z_39), .CK(clock), .Q(op_writeData[39])
         );
  DFF_X1 op_writeData_reg_231_ ( .D(n78), .CK(clock), .Q(op_writeData[231]) );
  DFF_X1 op_writeData_reg_167_ ( .D(U62_Z_167), .CK(clock), .Q(
        op_writeData[167]) );
  DFF_X1 op_writeData_reg_103_ ( .D(U62_Z_103), .CK(clock), .Q(
        op_writeData[103]) );
  DFF_X2 tempComputedDiagVal2_reg_38_ ( .D(n1266), .CK(clock), .QN(n404) );
  DFF_X1 op_writeData_reg_38_ ( .D(U62_Z_38), .CK(clock), .Q(op_writeData[38])
         );
  DFF_X1 op_writeData_reg_230_ ( .D(n77), .CK(clock), .Q(op_writeData[230]) );
  DFF_X1 op_writeData_reg_166_ ( .D(U62_Z_166), .CK(clock), .Q(
        op_writeData[166]) );
  DFF_X1 op_writeData_reg_102_ ( .D(U62_Z_102), .CK(clock), .Q(
        op_writeData[102]) );
  DFF_X2 tempComputedDiagVal2_reg_37_ ( .D(n1265), .CK(clock), .QN(n405) );
  DFF_X1 op_writeData_reg_37_ ( .D(U62_Z_37), .CK(clock), .Q(op_writeData[37])
         );
  DFF_X1 op_writeData_reg_229_ ( .D(n76), .CK(clock), .Q(op_writeData[229]) );
  DFF_X1 op_writeData_reg_165_ ( .D(U62_Z_165), .CK(clock), .Q(
        op_writeData[165]) );
  DFF_X1 op_writeData_reg_101_ ( .D(U62_Z_101), .CK(clock), .Q(
        op_writeData[101]) );
  DFF_X2 tempComputedDiagVal2_reg_36_ ( .D(n1264), .CK(clock), .QN(n406) );
  DFF_X1 op_writeData_reg_36_ ( .D(U62_Z_36), .CK(clock), .Q(op_writeData[36])
         );
  DFF_X1 op_writeData_reg_228_ ( .D(n75), .CK(clock), .Q(op_writeData[228]) );
  DFF_X1 op_writeData_reg_164_ ( .D(U62_Z_164), .CK(clock), .Q(
        op_writeData[164]) );
  DFF_X1 op_writeData_reg_100_ ( .D(U62_Z_100), .CK(clock), .Q(
        op_writeData[100]) );
  DFF_X2 tempComputedDiagVal2_reg_35_ ( .D(n1263), .CK(clock), .QN(n407) );
  DFF_X1 op_writeData_reg_99_ ( .D(U62_Z_99), .CK(clock), .Q(op_writeData[99])
         );
  DFF_X1 op_writeData_reg_35_ ( .D(U62_Z_35), .CK(clock), .Q(op_writeData[35])
         );
  DFF_X1 op_writeData_reg_227_ ( .D(n74), .CK(clock), .Q(op_writeData[227]) );
  DFF_X1 op_writeData_reg_163_ ( .D(U62_Z_163), .CK(clock), .Q(
        op_writeData[163]) );
  DFF_X2 tempComputedDiagVal2_reg_34_ ( .D(n1262), .CK(clock), .QN(n408) );
  DFF_X1 op_writeData_reg_98_ ( .D(U62_Z_98), .CK(clock), .Q(op_writeData[98])
         );
  DFF_X1 op_writeData_reg_34_ ( .D(U62_Z_34), .CK(clock), .Q(op_writeData[34])
         );
  DFF_X1 op_writeData_reg_226_ ( .D(n73), .CK(clock), .Q(op_writeData[226]) );
  DFF_X1 op_writeData_reg_162_ ( .D(U62_Z_162), .CK(clock), .Q(
        op_writeData[162]) );
  DFF_X2 tempComputedDiagVal2_reg_33_ ( .D(n1261), .CK(clock), .QN(n409) );
  DFF_X1 op_writeData_reg_97_ ( .D(U62_Z_97), .CK(clock), .Q(op_writeData[97])
         );
  DFF_X1 op_writeData_reg_33_ ( .D(U62_Z_33), .CK(clock), .Q(op_writeData[33])
         );
  DFF_X1 op_writeData_reg_225_ ( .D(n72), .CK(clock), .Q(op_writeData[225]) );
  DFF_X1 op_writeData_reg_161_ ( .D(U62_Z_161), .CK(clock), .Q(
        op_writeData[161]) );
  DFF_X2 tempComputedDiagVal2_reg_32_ ( .D(n1260), .CK(clock), .QN(n410) );
  DFF_X1 op_writeData_reg_96_ ( .D(U62_Z_96), .CK(clock), .Q(op_writeData[96])
         );
  DFF_X1 op_writeData_reg_32_ ( .D(U62_Z_32), .CK(clock), .Q(op_writeData[32])
         );
  DFF_X1 op_writeData_reg_224_ ( .D(n71), .CK(clock), .Q(op_writeData[224]) );
  DFF_X1 op_writeData_reg_160_ ( .D(U62_Z_160), .CK(clock), .Q(
        op_writeData[160]) );
  DFF_X2 tempComputedDiagVal2_reg_31_ ( .D(n1259), .CK(clock), .QN(n411) );
  DFF_X1 op_writeData_reg_95_ ( .D(U62_Z_95), .CK(clock), .Q(op_writeData[95])
         );
  DFF_X1 op_writeData_reg_31_ ( .D(U62_Z_31), .CK(clock), .Q(op_writeData[31])
         );
  DFF_X1 op_writeData_reg_223_ ( .D(n70), .CK(clock), .Q(op_writeData[223]) );
  DFF_X1 op_writeData_reg_159_ ( .D(U62_Z_159), .CK(clock), .Q(
        op_writeData[159]) );
  DFF_X2 tempComputedDiagVal2_reg_30_ ( .D(n1258), .CK(clock), .QN(n412) );
  DFF_X1 op_writeData_reg_94_ ( .D(U62_Z_94), .CK(clock), .Q(op_writeData[94])
         );
  DFF_X1 op_writeData_reg_30_ ( .D(U62_Z_30), .CK(clock), .Q(op_writeData[30])
         );
  DFF_X1 op_writeData_reg_222_ ( .D(n69), .CK(clock), .Q(op_writeData[222]) );
  DFF_X1 op_writeData_reg_158_ ( .D(U62_Z_158), .CK(clock), .Q(
        op_writeData[158]) );
  DFF_X2 tempComputedDiagVal2_reg_29_ ( .D(n1257), .CK(clock), .QN(n413) );
  DFF_X1 op_writeData_reg_93_ ( .D(U62_Z_93), .CK(clock), .Q(op_writeData[93])
         );
  DFF_X1 op_writeData_reg_29_ ( .D(U62_Z_29), .CK(clock), .Q(op_writeData[29])
         );
  DFF_X1 op_writeData_reg_221_ ( .D(n68), .CK(clock), .Q(op_writeData[221]) );
  DFF_X1 op_writeData_reg_157_ ( .D(U62_Z_157), .CK(clock), .Q(
        op_writeData[157]) );
  DFF_X2 tempComputedDiagVal2_reg_28_ ( .D(n1256), .CK(clock), .QN(n414) );
  DFF_X1 op_writeData_reg_92_ ( .D(U62_Z_92), .CK(clock), .Q(op_writeData[92])
         );
  DFF_X1 op_writeData_reg_28_ ( .D(U62_Z_28), .CK(clock), .Q(op_writeData[28])
         );
  DFF_X1 op_writeData_reg_220_ ( .D(n67), .CK(clock), .Q(op_writeData[220]) );
  DFF_X1 op_writeData_reg_156_ ( .D(U62_Z_156), .CK(clock), .Q(
        op_writeData[156]) );
  DFF_X2 tempComputedDiagVal2_reg_27_ ( .D(n1255), .CK(clock), .QN(n415) );
  DFF_X1 op_writeData_reg_91_ ( .D(U62_Z_91), .CK(clock), .Q(op_writeData[91])
         );
  DFF_X1 op_writeData_reg_27_ ( .D(U62_Z_27), .CK(clock), .Q(op_writeData[27])
         );
  DFF_X1 op_writeData_reg_219_ ( .D(n66), .CK(clock), .Q(op_writeData[219]) );
  DFF_X1 op_writeData_reg_155_ ( .D(U62_Z_155), .CK(clock), .Q(
        op_writeData[155]) );
  DFF_X2 tempComputedDiagVal2_reg_26_ ( .D(n1254), .CK(clock), .QN(n416) );
  DFF_X1 op_writeData_reg_90_ ( .D(U62_Z_90), .CK(clock), .Q(op_writeData[90])
         );
  DFF_X1 op_writeData_reg_26_ ( .D(U62_Z_26), .CK(clock), .Q(op_writeData[26])
         );
  DFF_X1 op_writeData_reg_218_ ( .D(n65), .CK(clock), .Q(op_writeData[218]) );
  DFF_X1 op_writeData_reg_154_ ( .D(U62_Z_154), .CK(clock), .Q(
        op_writeData[154]) );
  DFF_X2 tempComputedDiagVal2_reg_25_ ( .D(n1253), .CK(clock), .QN(n417) );
  DFF_X1 op_writeData_reg_89_ ( .D(U62_Z_89), .CK(clock), .Q(op_writeData[89])
         );
  DFF_X1 op_writeData_reg_25_ ( .D(U62_Z_25), .CK(clock), .Q(op_writeData[25])
         );
  DFF_X1 op_writeData_reg_217_ ( .D(n64), .CK(clock), .Q(op_writeData[217]) );
  DFF_X1 op_writeData_reg_153_ ( .D(U62_Z_153), .CK(clock), .Q(
        op_writeData[153]) );
  DFF_X2 tempComputedDiagVal2_reg_24_ ( .D(n1252), .CK(clock), .QN(n418) );
  DFF_X1 op_writeData_reg_88_ ( .D(U62_Z_88), .CK(clock), .Q(op_writeData[88])
         );
  DFF_X1 op_writeData_reg_24_ ( .D(U62_Z_24), .CK(clock), .Q(op_writeData[24])
         );
  DFF_X1 op_writeData_reg_216_ ( .D(n63), .CK(clock), .Q(op_writeData[216]) );
  DFF_X1 op_writeData_reg_152_ ( .D(U62_Z_152), .CK(clock), .Q(
        op_writeData[152]) );
  DFF_X2 tempComputedDiagVal2_reg_23_ ( .D(n1251), .CK(clock), .QN(n419) );
  DFF_X1 op_writeData_reg_87_ ( .D(U62_Z_87), .CK(clock), .Q(op_writeData[87])
         );
  DFF_X1 op_writeData_reg_23_ ( .D(U62_Z_23), .CK(clock), .Q(op_writeData[23])
         );
  DFF_X1 op_writeData_reg_215_ ( .D(n62), .CK(clock), .Q(op_writeData[215]) );
  DFF_X1 op_writeData_reg_151_ ( .D(U62_Z_151), .CK(clock), .Q(
        op_writeData[151]) );
  DFF_X2 tempComputedDiagVal2_reg_22_ ( .D(n1250), .CK(clock), .QN(n420) );
  DFF_X1 op_writeData_reg_86_ ( .D(U62_Z_86), .CK(clock), .Q(op_writeData[86])
         );
  DFF_X1 op_writeData_reg_22_ ( .D(U62_Z_22), .CK(clock), .Q(op_writeData[22])
         );
  DFF_X1 op_writeData_reg_214_ ( .D(n61), .CK(clock), .Q(op_writeData[214]) );
  DFF_X1 op_writeData_reg_150_ ( .D(U62_Z_150), .CK(clock), .Q(
        op_writeData[150]) );
  DFF_X2 tempComputedDiagVal2_reg_21_ ( .D(n1249), .CK(clock), .QN(n421) );
  DFF_X1 op_writeData_reg_85_ ( .D(U62_Z_85), .CK(clock), .Q(op_writeData[85])
         );
  DFF_X1 op_writeData_reg_213_ ( .D(n60), .CK(clock), .Q(op_writeData[213]) );
  DFF_X1 op_writeData_reg_21_ ( .D(U62_Z_21), .CK(clock), .Q(op_writeData[21])
         );
  DFF_X1 op_writeData_reg_149_ ( .D(U62_Z_149), .CK(clock), .Q(
        op_writeData[149]) );
  DFF_X2 tempComputedDiagVal2_reg_20_ ( .D(n1248), .CK(clock), .QN(n422) );
  DFF_X1 op_writeData_reg_84_ ( .D(U62_Z_84), .CK(clock), .Q(op_writeData[84])
         );
  DFF_X1 op_writeData_reg_212_ ( .D(n59), .CK(clock), .Q(op_writeData[212]) );
  DFF_X1 op_writeData_reg_20_ ( .D(U62_Z_20), .CK(clock), .Q(op_writeData[20])
         );
  DFF_X1 op_writeData_reg_148_ ( .D(U62_Z_148), .CK(clock), .Q(
        op_writeData[148]) );
  DFF_X2 tempComputedDiagVal2_reg_19_ ( .D(n1247), .CK(clock), .QN(n423) );
  DFF_X1 op_writeData_reg_83_ ( .D(U62_Z_83), .CK(clock), .Q(op_writeData[83])
         );
  DFF_X1 op_writeData_reg_211_ ( .D(n58), .CK(clock), .Q(op_writeData[211]) );
  DFF_X1 op_writeData_reg_19_ ( .D(U62_Z_19), .CK(clock), .Q(op_writeData[19])
         );
  DFF_X1 op_writeData_reg_147_ ( .D(U62_Z_147), .CK(clock), .Q(
        op_writeData[147]) );
  DFF_X2 tempComputedDiagVal2_reg_18_ ( .D(n1246), .CK(clock), .QN(n424) );
  DFF_X1 op_writeData_reg_82_ ( .D(U62_Z_82), .CK(clock), .Q(op_writeData[82])
         );
  DFF_X1 op_writeData_reg_210_ ( .D(n57), .CK(clock), .Q(op_writeData[210]) );
  DFF_X1 op_writeData_reg_18_ ( .D(U62_Z_18), .CK(clock), .Q(op_writeData[18])
         );
  DFF_X1 op_writeData_reg_146_ ( .D(U62_Z_146), .CK(clock), .Q(
        op_writeData[146]) );
  DFF_X2 tempComputedDiagVal2_reg_17_ ( .D(n1245), .CK(clock), .QN(n425) );
  DFF_X1 op_writeData_reg_81_ ( .D(U62_Z_81), .CK(clock), .Q(op_writeData[81])
         );
  DFF_X1 op_writeData_reg_209_ ( .D(n56), .CK(clock), .Q(op_writeData[209]) );
  DFF_X1 op_writeData_reg_17_ ( .D(U62_Z_17), .CK(clock), .Q(op_writeData[17])
         );
  DFF_X1 op_writeData_reg_145_ ( .D(U62_Z_145), .CK(clock), .Q(
        op_writeData[145]) );
  DFF_X2 tempComputedDiagVal2_reg_16_ ( .D(n1244), .CK(clock), .QN(n426) );
  DFF_X1 op_writeData_reg_80_ ( .D(U62_Z_80), .CK(clock), .Q(op_writeData[80])
         );
  DFF_X1 op_writeData_reg_208_ ( .D(n55), .CK(clock), .Q(op_writeData[208]) );
  DFF_X1 op_writeData_reg_16_ ( .D(U62_Z_16), .CK(clock), .Q(op_writeData[16])
         );
  DFF_X1 op_writeData_reg_144_ ( .D(U62_Z_144), .CK(clock), .Q(
        op_writeData[144]) );
  DFF_X2 tempComputedDiagVal2_reg_15_ ( .D(n1243), .CK(clock), .QN(n427) );
  DFF_X1 op_writeData_reg_79_ ( .D(U62_Z_79), .CK(clock), .Q(op_writeData[79])
         );
  DFF_X1 op_writeData_reg_207_ ( .D(n54), .CK(clock), .Q(op_writeData[207]) );
  DFF_X1 op_writeData_reg_15_ ( .D(U62_Z_15), .CK(clock), .Q(op_writeData[15])
         );
  DFF_X1 op_writeData_reg_143_ ( .D(U62_Z_143), .CK(clock), .Q(
        op_writeData[143]) );
  DFF_X2 tempComputedDiagVal2_reg_14_ ( .D(n1242), .CK(clock), .QN(n428) );
  DFF_X1 op_writeData_reg_78_ ( .D(U62_Z_78), .CK(clock), .Q(op_writeData[78])
         );
  DFF_X1 op_writeData_reg_206_ ( .D(n53), .CK(clock), .Q(op_writeData[206]) );
  DFF_X1 op_writeData_reg_142_ ( .D(U62_Z_142), .CK(clock), .Q(
        op_writeData[142]) );
  DFF_X1 op_writeData_reg_14_ ( .D(U62_Z_14), .CK(clock), .Q(op_writeData[14])
         );
  DFF_X2 tempComputedDiagVal2_reg_13_ ( .D(n1241), .CK(clock), .QN(n429) );
  DFF_X1 op_writeData_reg_77_ ( .D(U62_Z_77), .CK(clock), .Q(op_writeData[77])
         );
  DFF_X1 op_writeData_reg_205_ ( .D(n52), .CK(clock), .Q(op_writeData[205]) );
  DFF_X1 op_writeData_reg_141_ ( .D(U62_Z_141), .CK(clock), .Q(
        op_writeData[141]) );
  DFF_X1 op_writeData_reg_13_ ( .D(U62_Z_13), .CK(clock), .Q(op_writeData[13])
         );
  DFF_X2 tempComputedDiagVal2_reg_12_ ( .D(n1240), .CK(clock), .QN(n430) );
  DFF_X1 op_writeData_reg_76_ ( .D(U62_Z_76), .CK(clock), .Q(op_writeData[76])
         );
  DFF_X1 op_writeData_reg_204_ ( .D(n51), .CK(clock), .Q(op_writeData[204]) );
  DFF_X1 op_writeData_reg_140_ ( .D(U62_Z_140), .CK(clock), .Q(
        op_writeData[140]) );
  DFF_X1 op_writeData_reg_12_ ( .D(U62_Z_12), .CK(clock), .Q(op_writeData[12])
         );
  DFF_X2 tempComputedDiagVal2_reg_11_ ( .D(n1239), .CK(clock), .QN(n431) );
  DFF_X1 op_writeData_reg_75_ ( .D(U62_Z_75), .CK(clock), .Q(op_writeData[75])
         );
  DFF_X1 op_writeData_reg_203_ ( .D(n50), .CK(clock), .Q(op_writeData[203]) );
  DFF_X1 op_writeData_reg_139_ ( .D(U62_Z_139), .CK(clock), .Q(
        op_writeData[139]) );
  DFF_X1 op_writeData_reg_11_ ( .D(U62_Z_11), .CK(clock), .Q(op_writeData[11])
         );
  DFF_X2 tempComputedDiagVal2_reg_10_ ( .D(n1238), .CK(clock), .QN(n432) );
  DFF_X1 op_writeData_reg_74_ ( .D(U62_Z_74), .CK(clock), .Q(op_writeData[74])
         );
  DFF_X1 op_writeData_reg_202_ ( .D(n49), .CK(clock), .Q(op_writeData[202]) );
  DFF_X1 op_writeData_reg_138_ ( .D(U62_Z_138), .CK(clock), .Q(
        op_writeData[138]) );
  DFF_X1 op_writeData_reg_10_ ( .D(U62_Z_10), .CK(clock), .Q(op_writeData[10])
         );
  DFF_X2 tempComputedDiagVal2_reg_9_ ( .D(n1237), .CK(clock), .QN(n433) );
  DFF_X1 op_writeData_reg_9_ ( .D(U62_Z_9), .CK(clock), .Q(op_writeData[9]) );
  DFF_X1 op_writeData_reg_73_ ( .D(U62_Z_73), .CK(clock), .Q(op_writeData[73])
         );
  DFF_X1 op_writeData_reg_201_ ( .D(n48), .CK(clock), .Q(op_writeData[201]) );
  DFF_X1 op_writeData_reg_137_ ( .D(U62_Z_137), .CK(clock), .Q(
        op_writeData[137]) );
  DFF_X2 tempComputedDiagVal2_reg_8_ ( .D(n1236), .CK(clock), .QN(n434) );
  DFF_X1 op_writeData_reg_8_ ( .D(U62_Z_8), .CK(clock), .Q(op_writeData[8]) );
  DFF_X1 op_writeData_reg_72_ ( .D(U62_Z_72), .CK(clock), .Q(op_writeData[72])
         );
  DFF_X1 op_writeData_reg_200_ ( .D(n47), .CK(clock), .Q(op_writeData[200]) );
  DFF_X1 op_writeData_reg_136_ ( .D(U62_Z_136), .CK(clock), .Q(
        op_writeData[136]) );
  DFF_X2 tempComputedDiagVal2_reg_7_ ( .D(n1235), .CK(clock), .QN(n435) );
  DFF_X1 op_writeData_reg_71_ ( .D(U62_Z_71), .CK(clock), .Q(op_writeData[71])
         );
  DFF_X1 op_writeData_reg_7_ ( .D(U62_Z_7), .CK(clock), .Q(op_writeData[7]) );
  DFF_X1 op_writeData_reg_199_ ( .D(n46), .CK(clock), .Q(op_writeData[199]) );
  DFF_X1 op_writeData_reg_135_ ( .D(U62_Z_135), .CK(clock), .Q(
        op_writeData[135]) );
  DFF_X2 tempComputedDiagVal2_reg_6_ ( .D(n1234), .CK(clock), .QN(n436) );
  DFF_X1 op_writeData_reg_70_ ( .D(U62_Z_70), .CK(clock), .Q(op_writeData[70])
         );
  DFF_X1 op_writeData_reg_6_ ( .D(U62_Z_6), .CK(clock), .Q(op_writeData[6]) );
  DFF_X1 op_writeData_reg_198_ ( .D(n45), .CK(clock), .Q(op_writeData[198]) );
  DFF_X1 op_writeData_reg_134_ ( .D(U62_Z_134), .CK(clock), .Q(
        op_writeData[134]) );
  DFF_X2 tempComputedDiagVal2_reg_5_ ( .D(n1233), .CK(clock), .QN(n437) );
  DFF_X1 op_writeData_reg_69_ ( .D(U62_Z_69), .CK(clock), .Q(op_writeData[69])
         );
  DFF_X1 op_writeData_reg_5_ ( .D(U62_Z_5), .CK(clock), .Q(op_writeData[5]) );
  DFF_X1 op_writeData_reg_197_ ( .D(n44), .CK(clock), .Q(op_writeData[197]) );
  DFF_X1 op_writeData_reg_133_ ( .D(U62_Z_133), .CK(clock), .Q(
        op_writeData[133]) );
  DFF_X2 tempComputedDiagVal2_reg_4_ ( .D(n1232), .CK(clock), .QN(n438) );
  DFF_X1 op_writeData_reg_68_ ( .D(U62_Z_68), .CK(clock), .Q(op_writeData[68])
         );
  DFF_X1 op_writeData_reg_4_ ( .D(U62_Z_4), .CK(clock), .Q(op_writeData[4]) );
  DFF_X1 op_writeData_reg_196_ ( .D(n43), .CK(clock), .Q(op_writeData[196]) );
  DFF_X1 op_writeData_reg_132_ ( .D(U62_Z_132), .CK(clock), .Q(
        op_writeData[132]) );
  DFF_X2 tempComputedDiagVal2_reg_3_ ( .D(n1231), .CK(clock), .QN(n439) );
  DFF_X1 op_writeData_reg_67_ ( .D(U62_Z_67), .CK(clock), .Q(op_writeData[67])
         );
  DFF_X1 op_writeData_reg_3_ ( .D(U62_Z_3), .CK(clock), .Q(op_writeData[3]) );
  DFF_X1 op_writeData_reg_195_ ( .D(n42), .CK(clock), .Q(op_writeData[195]) );
  DFF_X1 op_writeData_reg_131_ ( .D(U62_Z_131), .CK(clock), .Q(
        op_writeData[131]) );
  DFF_X2 tempComputedDiagVal2_reg_2_ ( .D(n1230), .CK(clock), .QN(n440) );
  DFF_X1 op_writeData_reg_66_ ( .D(U62_Z_66), .CK(clock), .Q(op_writeData[66])
         );
  DFF_X1 op_writeData_reg_2_ ( .D(U62_Z_2), .CK(clock), .Q(op_writeData[2]) );
  DFF_X1 op_writeData_reg_194_ ( .D(n41), .CK(clock), .Q(op_writeData[194]) );
  DFF_X1 op_writeData_reg_130_ ( .D(U62_Z_130), .CK(clock), .Q(
        op_writeData[130]) );
  DFF_X2 tempComputedDiagVal2_reg_1_ ( .D(n1229), .CK(clock), .QN(n441) );
  DFF_X1 op_writeData_reg_65_ ( .D(U62_Z_65), .CK(clock), .Q(op_writeData[65])
         );
  DFF_X1 op_writeData_reg_193_ ( .D(n40), .CK(clock), .Q(op_writeData[193]) );
  DFF_X1 op_writeData_reg_129_ ( .D(U62_Z_129), .CK(clock), .Q(
        op_writeData[129]) );
  DFF_X1 op_writeData_reg_1_ ( .D(U62_Z_1), .CK(clock), .Q(op_writeData[1]) );
  DFF_X2 tempComputedDiagVal2_reg_0_ ( .D(n1228), .CK(clock), .QN(n442) );
  DFF_X1 op_writeData_reg_64_ ( .D(U62_Z_64), .CK(clock), .Q(op_writeData[64])
         );
  DFF_X1 op_writeData_reg_192_ ( .D(n39), .CK(clock), .Q(op_writeData[192]) );
  DFF_X1 op_writeData_reg_128_ ( .D(U62_Z_128), .CK(clock), .Q(
        op_writeData[128]) );
  DFF_X1 op_writeData_reg_0_ ( .D(U62_Z_0), .CK(clock), .Q(op_writeData[0]) );
  OAI22_X2 U6 ( .A1(n4315), .A2(n442), .B1(n4313), .B2(n716), .ZN(n1228) );
  OAI22_X2 U7 ( .A1(n765), .A2(n441), .B1(n4312), .B2(n715), .ZN(n1229) );
  OAI22_X2 U8 ( .A1(n765), .A2(n440), .B1(n4313), .B2(n714), .ZN(n1230) );
  OAI22_X2 U9 ( .A1(n765), .A2(n439), .B1(n4312), .B2(n713), .ZN(n1231) );
  OAI22_X2 U10 ( .A1(n765), .A2(n438), .B1(n4313), .B2(n712), .ZN(n1232) );
  OAI22_X2 U11 ( .A1(n4315), .A2(n437), .B1(n4313), .B2(n711), .ZN(n1233) );
  OAI22_X2 U12 ( .A1(n4314), .A2(n436), .B1(n4313), .B2(n710), .ZN(n1234) );
  OAI22_X2 U13 ( .A1(n4315), .A2(n435), .B1(n4312), .B2(n709), .ZN(n1235) );
  OAI22_X2 U14 ( .A1(n4315), .A2(n434), .B1(n4313), .B2(n708), .ZN(n1236) );
  OAI22_X2 U15 ( .A1(n4314), .A2(n433), .B1(n4313), .B2(n707), .ZN(n1237) );
  OAI22_X2 U16 ( .A1(n4315), .A2(n432), .B1(n4313), .B2(n706), .ZN(n1238) );
  OAI22_X2 U17 ( .A1(n4314), .A2(n431), .B1(n4313), .B2(n705), .ZN(n1239) );
  OAI22_X2 U18 ( .A1(n4315), .A2(n430), .B1(n4313), .B2(n704), .ZN(n1240) );
  OAI22_X2 U19 ( .A1(n4314), .A2(n429), .B1(n4313), .B2(n703), .ZN(n1241) );
  OAI22_X2 U20 ( .A1(n4315), .A2(n428), .B1(n4313), .B2(n702), .ZN(n1242) );
  OAI22_X2 U21 ( .A1(n4314), .A2(n427), .B1(n4313), .B2(n701), .ZN(n1243) );
  OAI22_X2 U22 ( .A1(n4315), .A2(n426), .B1(n4313), .B2(n700), .ZN(n1244) );
  OAI22_X2 U23 ( .A1(n4314), .A2(n425), .B1(n4313), .B2(n699), .ZN(n1245) );
  OAI22_X2 U24 ( .A1(n4314), .A2(n424), .B1(n4313), .B2(n698), .ZN(n1246) );
  OAI22_X2 U25 ( .A1(n4315), .A2(n423), .B1(n4313), .B2(n697), .ZN(n1247) );
  OAI22_X2 U26 ( .A1(n4314), .A2(n422), .B1(n4313), .B2(n696), .ZN(n1248) );
  OAI22_X2 U27 ( .A1(n4315), .A2(n421), .B1(n4313), .B2(n695), .ZN(n1249) );
  OAI22_X2 U28 ( .A1(n4314), .A2(n420), .B1(n4313), .B2(n694), .ZN(n1250) );
  OAI22_X2 U29 ( .A1(n4315), .A2(n419), .B1(n4313), .B2(n693), .ZN(n1251) );
  OAI22_X2 U30 ( .A1(n4314), .A2(n418), .B1(n4313), .B2(n692), .ZN(n1252) );
  OAI22_X2 U31 ( .A1(n4315), .A2(n417), .B1(n4312), .B2(n691), .ZN(n1253) );
  OAI22_X2 U32 ( .A1(n4315), .A2(n416), .B1(n4313), .B2(n690), .ZN(n1254) );
  OAI22_X2 U33 ( .A1(n4314), .A2(n415), .B1(n4312), .B2(n689), .ZN(n1255) );
  OAI22_X2 U34 ( .A1(n4315), .A2(n414), .B1(n4312), .B2(n688), .ZN(n1256) );
  OAI22_X2 U35 ( .A1(n4314), .A2(n413), .B1(n4313), .B2(n687), .ZN(n1257) );
  OAI22_X2 U36 ( .A1(n4315), .A2(n412), .B1(n4313), .B2(n686), .ZN(n1258) );
  OAI22_X2 U37 ( .A1(n4314), .A2(n411), .B1(n4312), .B2(n685), .ZN(n1259) );
  OAI22_X2 U38 ( .A1(n4315), .A2(n410), .B1(n4313), .B2(n684), .ZN(n1260) );
  OAI22_X2 U39 ( .A1(n4314), .A2(n409), .B1(n4312), .B2(n683), .ZN(n1261) );
  OAI22_X2 U40 ( .A1(n4315), .A2(n408), .B1(n4312), .B2(n682), .ZN(n1262) );
  OAI22_X2 U41 ( .A1(n4314), .A2(n407), .B1(n4313), .B2(n681), .ZN(n1263) );
  OAI22_X2 U42 ( .A1(n4315), .A2(n406), .B1(n4313), .B2(n680), .ZN(n1264) );
  OAI22_X2 U43 ( .A1(n4314), .A2(n405), .B1(n4312), .B2(n679), .ZN(n1265) );
  OAI22_X2 U44 ( .A1(n4314), .A2(n404), .B1(n4313), .B2(n678), .ZN(n1266) );
  OAI22_X2 U45 ( .A1(n4315), .A2(n403), .B1(n4312), .B2(n677), .ZN(n1267) );
  OAI22_X2 U46 ( .A1(n4315), .A2(n402), .B1(n4313), .B2(n676), .ZN(n1268) );
  OAI22_X2 U47 ( .A1(n4314), .A2(n401), .B1(n4312), .B2(n675), .ZN(n1269) );
  OAI22_X2 U48 ( .A1(n4314), .A2(n400), .B1(n4313), .B2(n674), .ZN(n1270) );
  OAI22_X2 U49 ( .A1(n4315), .A2(n399), .B1(n4312), .B2(n673), .ZN(n1271) );
  OAI22_X2 U50 ( .A1(n4314), .A2(n398), .B1(n4313), .B2(n672), .ZN(n1272) );
  OAI22_X2 U51 ( .A1(n4314), .A2(n397), .B1(n4312), .B2(n671), .ZN(n1273) );
  OAI22_X2 U52 ( .A1(n4315), .A2(n396), .B1(n4313), .B2(n670), .ZN(n1274) );
  OAI22_X2 U53 ( .A1(n4315), .A2(n395), .B1(n4312), .B2(n669), .ZN(n1275) );
  OAI22_X2 U54 ( .A1(n4310), .A2(n394), .B1(n716), .B2(n4308), .ZN(n1276) );
  OAI22_X2 U55 ( .A1(n4311), .A2(n393), .B1(n715), .B2(n4309), .ZN(n1277) );
  OAI22_X2 U56 ( .A1(n4311), .A2(n392), .B1(n714), .B2(n4308), .ZN(n1278) );
  OAI22_X2 U57 ( .A1(n4311), .A2(n391), .B1(n713), .B2(n4308), .ZN(n1279) );
  OAI22_X2 U58 ( .A1(n4311), .A2(n390), .B1(n712), .B2(n4309), .ZN(n1280) );
  OAI22_X2 U59 ( .A1(n4310), .A2(n389), .B1(n711), .B2(n4308), .ZN(n1281) );
  OAI22_X2 U60 ( .A1(n4311), .A2(n388), .B1(n710), .B2(n4308), .ZN(n1282) );
  OAI22_X2 U61 ( .A1(n4310), .A2(n387), .B1(n709), .B2(n4309), .ZN(n1283) );
  OAI22_X2 U62 ( .A1(n4311), .A2(n386), .B1(n708), .B2(n4308), .ZN(n1284) );
  OAI22_X2 U63 ( .A1(n4310), .A2(n385), .B1(n707), .B2(n4309), .ZN(n1285) );
  OAI22_X2 U64 ( .A1(n4310), .A2(n384), .B1(n706), .B2(n4309), .ZN(n1286) );
  OAI22_X2 U65 ( .A1(n4311), .A2(n383), .B1(n705), .B2(n4308), .ZN(n1287) );
  OAI22_X2 U66 ( .A1(n4311), .A2(n382), .B1(n704), .B2(n4308), .ZN(n1288) );
  OAI22_X2 U67 ( .A1(n4311), .A2(n381), .B1(n703), .B2(n4309), .ZN(n1289) );
  OAI22_X2 U68 ( .A1(n4311), .A2(n380), .B1(n702), .B2(n4308), .ZN(n1290) );
  OAI22_X2 U69 ( .A1(n4311), .A2(n379), .B1(n701), .B2(n4309), .ZN(n1291) );
  OAI22_X2 U70 ( .A1(n4311), .A2(n378), .B1(n700), .B2(n4309), .ZN(n1292) );
  OAI22_X2 U71 ( .A1(n4311), .A2(n377), .B1(n699), .B2(n4308), .ZN(n1293) );
  OAI22_X2 U72 ( .A1(n4311), .A2(n376), .B1(n698), .B2(n4308), .ZN(n1294) );
  OAI22_X2 U73 ( .A1(n4311), .A2(n375), .B1(n697), .B2(n4309), .ZN(n1295) );
  OAI22_X2 U74 ( .A1(n4311), .A2(n374), .B1(n696), .B2(n4309), .ZN(n1296) );
  OAI22_X2 U75 ( .A1(n4311), .A2(n373), .B1(n695), .B2(n4309), .ZN(n1297) );
  OAI22_X2 U76 ( .A1(n4311), .A2(n372), .B1(n694), .B2(n4308), .ZN(n1298) );
  OAI22_X2 U77 ( .A1(n4311), .A2(n371), .B1(n693), .B2(n4309), .ZN(n1299) );
  OAI22_X2 U78 ( .A1(n4310), .A2(n370), .B1(n692), .B2(n4308), .ZN(n1300) );
  OAI22_X2 U79 ( .A1(n4310), .A2(n369), .B1(n691), .B2(n4308), .ZN(n1301) );
  OAI22_X2 U80 ( .A1(n4310), .A2(n368), .B1(n690), .B2(n4308), .ZN(n1302) );
  OAI22_X2 U81 ( .A1(n4310), .A2(n367), .B1(n689), .B2(n4308), .ZN(n1303) );
  OAI22_X2 U82 ( .A1(n4310), .A2(n366), .B1(n688), .B2(n4308), .ZN(n1304) );
  OAI22_X2 U83 ( .A1(n4310), .A2(n365), .B1(n687), .B2(n4308), .ZN(n1305) );
  OAI22_X2 U84 ( .A1(n4310), .A2(n364), .B1(n686), .B2(n4308), .ZN(n1306) );
  OAI22_X2 U85 ( .A1(n4310), .A2(n363), .B1(n685), .B2(n4308), .ZN(n1307) );
  OAI22_X2 U86 ( .A1(n4310), .A2(n362), .B1(n684), .B2(n4308), .ZN(n1308) );
  OAI22_X2 U87 ( .A1(n4310), .A2(n361), .B1(n683), .B2(n4308), .ZN(n1309) );
  OAI22_X2 U88 ( .A1(n4310), .A2(n360), .B1(n682), .B2(n4308), .ZN(n1310) );
  OAI22_X2 U89 ( .A1(n4310), .A2(n359), .B1(n681), .B2(n4308), .ZN(n1311) );
  OAI22_X2 U90 ( .A1(n4311), .A2(n358), .B1(n680), .B2(n4309), .ZN(n1312) );
  OAI22_X2 U91 ( .A1(n4310), .A2(n357), .B1(n679), .B2(n4309), .ZN(n1313) );
  OAI22_X2 U92 ( .A1(n4311), .A2(n356), .B1(n678), .B2(n4309), .ZN(n1314) );
  OAI22_X2 U93 ( .A1(n4311), .A2(n355), .B1(n677), .B2(n4309), .ZN(n1315) );
  OAI22_X2 U94 ( .A1(n4310), .A2(n354), .B1(n676), .B2(n4309), .ZN(n1316) );
  OAI22_X2 U95 ( .A1(n4310), .A2(n353), .B1(n675), .B2(n4309), .ZN(n1317) );
  OAI22_X2 U96 ( .A1(n4311), .A2(n352), .B1(n674), .B2(n4309), .ZN(n1318) );
  OAI22_X2 U97 ( .A1(n4310), .A2(n351), .B1(n673), .B2(n4309), .ZN(n1319) );
  OAI22_X2 U98 ( .A1(n4311), .A2(n350), .B1(n672), .B2(n4309), .ZN(n1320) );
  OAI22_X2 U99 ( .A1(n4311), .A2(n349), .B1(n671), .B2(n4309), .ZN(n1321) );
  OAI22_X2 U100 ( .A1(n4310), .A2(n348), .B1(n670), .B2(n4309), .ZN(n1322) );
  OAI22_X2 U101 ( .A1(n4310), .A2(n347), .B1(n669), .B2(n4309), .ZN(n1323) );
  OAI22_X2 U102 ( .A1(n4314), .A2(n346), .B1(n4313), .B2(n476), .ZN(n1324) );
  OAI22_X2 U103 ( .A1(n4314), .A2(n345), .B1(n4312), .B2(n475), .ZN(n1325) );
  OAI22_X2 U104 ( .A1(n4315), .A2(n344), .B1(n4313), .B2(n474), .ZN(n1326) );
  OAI22_X2 U105 ( .A1(n4315), .A2(n343), .B1(n4312), .B2(n473), .ZN(n1327) );
  OAI22_X2 U106 ( .A1(n4311), .A2(n342), .B1(n4309), .B2(n476), .ZN(n1328) );
  OAI22_X2 U107 ( .A1(n4310), .A2(n341), .B1(n4308), .B2(n475), .ZN(n1329) );
  OAI22_X2 U108 ( .A1(n4311), .A2(n340), .B1(n4309), .B2(n474), .ZN(n1330) );
  OAI22_X2 U109 ( .A1(n4310), .A2(n339), .B1(n4309), .B2(n473), .ZN(n1331) );
  OAI22_X2 U110 ( .A1(n4314), .A2(n338), .B1(n4313), .B2(n472), .ZN(n1332) );
  OAI22_X2 U111 ( .A1(n4314), .A2(n337), .B1(n4312), .B2(n471), .ZN(n1333) );
  OAI22_X2 U112 ( .A1(n4315), .A2(n336), .B1(n4312), .B2(n470), .ZN(n1334) );
  OAI22_X2 U113 ( .A1(n4314), .A2(n335), .B1(n4312), .B2(n469), .ZN(n1335) );
  OAI22_X2 U114 ( .A1(n4311), .A2(n334), .B1(n4308), .B2(n472), .ZN(n1336) );
  OAI22_X2 U115 ( .A1(n4310), .A2(n333), .B1(n4308), .B2(n471), .ZN(n1337) );
  OAI22_X2 U116 ( .A1(n4311), .A2(n332), .B1(n4309), .B2(n470), .ZN(n1338) );
  OAI22_X2 U117 ( .A1(n4310), .A2(n331), .B1(n4308), .B2(n469), .ZN(n1339) );
  OAI221_X2 U118 ( .B1(n4312), .B2(n467), .C1(n4315), .C2(n329), .A(n769), 
        .ZN(n1340) );
  OAI221_X2 U119 ( .B1(n4312), .B2(n466), .C1(n4314), .C2(n328), .A(n4289), 
        .ZN(n1341) );
  OAI221_X2 U120 ( .B1(n4312), .B2(n465), .C1(n4315), .C2(n327), .A(n769), 
        .ZN(n1342) );
  OAI221_X2 U121 ( .B1(n4312), .B2(n464), .C1(n4314), .C2(n326), .A(n4289), 
        .ZN(n1343) );
  OAI221_X2 U122 ( .B1(n4312), .B2(n463), .C1(n4315), .C2(n325), .A(n769), 
        .ZN(n1344) );
  OAI221_X2 U123 ( .B1(n4312), .B2(n462), .C1(n4314), .C2(n324), .A(n4289), 
        .ZN(n1345) );
  OAI221_X2 U124 ( .B1(n4312), .B2(n461), .C1(n4315), .C2(n323), .A(n769), 
        .ZN(n1346) );
  OAI221_X2 U125 ( .B1(n4312), .B2(n460), .C1(n4314), .C2(n322), .A(n4289), 
        .ZN(n1347) );
  OAI221_X2 U126 ( .B1(n4312), .B2(n459), .C1(n4315), .C2(n321), .A(n769), 
        .ZN(n1348) );
  OAI221_X2 U127 ( .B1(n4312), .B2(n458), .C1(n4314), .C2(n320), .A(n4289), 
        .ZN(n1349) );
  OAI221_X2 U128 ( .B1(n4312), .B2(n457), .C1(n4315), .C2(n308), .A(n769), 
        .ZN(n1350) );
  OAI221_X2 U129 ( .B1(n4312), .B2(n456), .C1(n4314), .C2(n307), .A(n4289), 
        .ZN(n1351) );
  OAI221_X2 U130 ( .B1(n4312), .B2(n455), .C1(n4315), .C2(n306), .A(n769), 
        .ZN(n1352) );
  OAI221_X2 U131 ( .B1(n4313), .B2(n454), .C1(n4314), .C2(n305), .A(n4289), 
        .ZN(n1353) );
  OAI221_X2 U132 ( .B1(n4312), .B2(n453), .C1(n4314), .C2(n304), .A(n769), 
        .ZN(n1354) );
  OAI221_X2 U133 ( .B1(n4312), .B2(n452), .C1(n4315), .C2(n303), .A(n4289), 
        .ZN(n1355) );
  OAI221_X2 U134 ( .B1(n4313), .B2(n451), .C1(n4315), .C2(n302), .A(n769), 
        .ZN(n1356) );
  OAI221_X2 U135 ( .B1(n4313), .B2(n450), .C1(n4314), .C2(n301), .A(n4289), 
        .ZN(n1357) );
  OAI221_X2 U136 ( .B1(n4312), .B2(n449), .C1(n4314), .C2(n300), .A(n769), 
        .ZN(n1358) );
  OAI221_X2 U137 ( .B1(n4312), .B2(n448), .C1(n4315), .C2(n299), .A(n4289), 
        .ZN(n1359) );
  OAI221_X2 U138 ( .B1(n4312), .B2(n447), .C1(n4315), .C2(n298), .A(n769), 
        .ZN(n1360) );
  OAI22_X2 U139 ( .A1(n4311), .A2(n319), .B1(n4309), .B2(n468), .ZN(n1361) );
  OAI22_X2 U140 ( .A1(n4310), .A2(n318), .B1(n4309), .B2(n467), .ZN(n1362) );
  OAI22_X2 U141 ( .A1(n4311), .A2(n317), .B1(n4308), .B2(n466), .ZN(n1363) );
  OAI22_X2 U142 ( .A1(n4310), .A2(n316), .B1(n4308), .B2(n465), .ZN(n1364) );
  OAI22_X2 U143 ( .A1(n4311), .A2(n315), .B1(n4309), .B2(n464), .ZN(n1365) );
  OAI22_X2 U144 ( .A1(n4311), .A2(n314), .B1(n4308), .B2(n463), .ZN(n1366) );
  OAI22_X2 U145 ( .A1(n4311), .A2(n313), .B1(n4309), .B2(n462), .ZN(n1367) );
  OAI22_X2 U146 ( .A1(n4311), .A2(n312), .B1(n4308), .B2(n461), .ZN(n1368) );
  OAI22_X2 U147 ( .A1(n4311), .A2(n311), .B1(n4309), .B2(n460), .ZN(n1369) );
  OAI22_X2 U148 ( .A1(n4311), .A2(n310), .B1(n4308), .B2(n459), .ZN(n1370) );
  OAI22_X2 U149 ( .A1(n4311), .A2(n309), .B1(n4309), .B2(n458), .ZN(n1371) );
  OAI22_X2 U150 ( .A1(n4311), .A2(n297), .B1(n4308), .B2(n457), .ZN(n1372) );
  OAI22_X2 U151 ( .A1(n4311), .A2(n296), .B1(n4309), .B2(n456), .ZN(n1373) );
  OAI22_X2 U152 ( .A1(n4311), .A2(n295), .B1(n4308), .B2(n455), .ZN(n1374) );
  OAI22_X2 U153 ( .A1(n4311), .A2(n294), .B1(n4309), .B2(n454), .ZN(n1375) );
  OAI22_X2 U154 ( .A1(n4311), .A2(n293), .B1(n4308), .B2(n453), .ZN(n1376) );
  OAI22_X2 U155 ( .A1(n4310), .A2(n292), .B1(n4309), .B2(n452), .ZN(n1377) );
  OAI22_X2 U156 ( .A1(n4311), .A2(n291), .B1(n4308), .B2(n451), .ZN(n1378) );
  OAI22_X2 U157 ( .A1(n4311), .A2(n290), .B1(n4308), .B2(n450), .ZN(n1379) );
  OAI22_X2 U158 ( .A1(n4311), .A2(n289), .B1(n4309), .B2(n449), .ZN(n1380) );
  OAI22_X2 U159 ( .A1(n4310), .A2(n288), .B1(n4309), .B2(n448), .ZN(n1381) );
  OAI22_X2 U160 ( .A1(n4311), .A2(n287), .B1(n4308), .B2(n447), .ZN(n1382) );
  OAI22_X2 U164 ( .A1(n121), .A2(n4318), .B1(n4320), .B2(n774), .ZN(n1383) );
  OAI221_X2 U165 ( .B1(n4313), .B2(n468), .C1(n4314), .C2(n330), .A(n4289), 
        .ZN(n1384) );
  NAND3_X2 U166 ( .A1(n4315), .A2(reset), .A3(n771), .ZN(n769) );
  NOR3_X2 U169 ( .A1(n772), .A2(n771), .A3(n775), .ZN(n776) );
  NOR2_X2 U170 ( .A1(n446), .A2(n445), .ZN(n775) );
  NOR2_X2 U171 ( .A1(n446), .A2(cpDoneFlag), .ZN(n771) );
  NAND2_X2 U172 ( .A1(n777), .A2(n778), .ZN(n773) );
  OAI221_X2 U173 ( .B1(n4333), .B2(n729), .C1(n4297), .C2(n186), .A(n780), 
        .ZN(U62_Z_99) );
  OAI221_X2 U175 ( .B1(n4333), .B2(n730), .C1(n4297), .C2(n187), .A(n784), 
        .ZN(U62_Z_98) );
  OAI221_X2 U177 ( .B1(n4333), .B2(n731), .C1(n4297), .C2(n188), .A(n786), 
        .ZN(U62_Z_97) );
  OAI221_X2 U179 ( .B1(n4333), .B2(n732), .C1(n4297), .C2(n189), .A(n788), 
        .ZN(U62_Z_96) );
  OAI221_X2 U181 ( .B1(n4333), .B2(n733), .C1(n4297), .C2(n190), .A(n790), 
        .ZN(U62_Z_95) );
  OAI221_X2 U183 ( .B1(n4333), .B2(n734), .C1(n4297), .C2(n191), .A(n792), 
        .ZN(U62_Z_94) );
  OAI221_X2 U185 ( .B1(n4333), .B2(n735), .C1(n4297), .C2(n192), .A(n794), 
        .ZN(U62_Z_93) );
  OAI221_X2 U187 ( .B1(n4333), .B2(n736), .C1(n4297), .C2(n193), .A(n796), 
        .ZN(U62_Z_92) );
  OAI221_X2 U189 ( .B1(n4333), .B2(n737), .C1(n4297), .C2(n194), .A(n798), 
        .ZN(U62_Z_91) );
  OAI221_X2 U191 ( .B1(n4333), .B2(n738), .C1(n4297), .C2(n195), .A(n800), 
        .ZN(U62_Z_90) );
  OAI221_X2 U193 ( .B1(n4302), .B2(n755), .C1(n4297), .C2(n260), .A(n803), 
        .ZN(U62_Z_9) );
  OAI221_X2 U195 ( .B1(n4333), .B2(n739), .C1(n4299), .C2(n196), .A(n807), 
        .ZN(U62_Z_89) );
  OAI221_X2 U197 ( .B1(n4333), .B2(n740), .C1(n4297), .C2(n197), .A(n809), 
        .ZN(U62_Z_88) );
  OAI221_X2 U199 ( .B1(n4333), .B2(n741), .C1(n4297), .C2(n198), .A(n811), 
        .ZN(U62_Z_87) );
  OAI221_X2 U201 ( .B1(n4333), .B2(n742), .C1(n4298), .C2(n199), .A(n813), 
        .ZN(U62_Z_86) );
  OAI221_X2 U203 ( .B1(n4333), .B2(n743), .C1(n4297), .C2(n200), .A(n815), 
        .ZN(U62_Z_85) );
  OAI221_X2 U205 ( .B1(n4333), .B2(n744), .C1(n4298), .C2(n201), .A(n817), 
        .ZN(U62_Z_84) );
  OAI221_X2 U207 ( .B1(n4333), .B2(n745), .C1(n4298), .C2(n202), .A(n819), 
        .ZN(U62_Z_83) );
  OAI221_X2 U209 ( .B1(n4333), .B2(n746), .C1(n4297), .C2(n203), .A(n821), 
        .ZN(U62_Z_82) );
  OAI221_X2 U211 ( .B1(n4333), .B2(n747), .C1(n4297), .C2(n204), .A(n823), 
        .ZN(U62_Z_81) );
  OAI221_X2 U213 ( .B1(n4333), .B2(n748), .C1(n4298), .C2(n205), .A(n825), 
        .ZN(U62_Z_80) );
  OAI221_X2 U215 ( .B1(n4302), .B2(n756), .C1(n4297), .C2(n261), .A(n827), 
        .ZN(U62_Z_8) );
  OAI221_X2 U217 ( .B1(n4333), .B2(n749), .C1(n4297), .C2(n206), .A(n829), 
        .ZN(U62_Z_79) );
  OAI221_X2 U219 ( .B1(n4333), .B2(n750), .C1(n4297), .C2(n207), .A(n831), 
        .ZN(U62_Z_78) );
  OAI221_X2 U221 ( .B1(n4333), .B2(n751), .C1(n4297), .C2(n208), .A(n833), 
        .ZN(U62_Z_77) );
  OAI221_X2 U223 ( .B1(n4333), .B2(n752), .C1(n4298), .C2(n209), .A(n835), 
        .ZN(U62_Z_76) );
  OAI221_X2 U225 ( .B1(n4333), .B2(n753), .C1(n4298), .C2(n210), .A(n837), 
        .ZN(U62_Z_75) );
  OAI221_X2 U227 ( .B1(n4333), .B2(n754), .C1(n4298), .C2(n211), .A(n839), 
        .ZN(U62_Z_74) );
  OAI221_X2 U229 ( .B1(n4333), .B2(n755), .C1(n4298), .C2(n212), .A(n841), 
        .ZN(U62_Z_73) );
  OAI221_X2 U231 ( .B1(n4333), .B2(n756), .C1(n4298), .C2(n213), .A(n842), 
        .ZN(U62_Z_72) );
  OAI221_X2 U233 ( .B1(n4333), .B2(n757), .C1(n4298), .C2(n214), .A(n843), 
        .ZN(U62_Z_71) );
  OAI221_X2 U235 ( .B1(n4333), .B2(n758), .C1(n4298), .C2(n215), .A(n845), 
        .ZN(U62_Z_70) );
  OAI221_X2 U237 ( .B1(n4302), .B2(n757), .C1(n4298), .C2(n262), .A(n847), 
        .ZN(U62_Z_7) );
  OAI221_X2 U239 ( .B1(n4333), .B2(n759), .C1(n4298), .C2(n216), .A(n848), 
        .ZN(U62_Z_69) );
  OAI221_X2 U241 ( .B1(n4333), .B2(n760), .C1(n4298), .C2(n217), .A(n850), 
        .ZN(U62_Z_68) );
  OAI221_X2 U243 ( .B1(n4333), .B2(n761), .C1(n4298), .C2(n218), .A(n852), 
        .ZN(U62_Z_67) );
  OAI221_X2 U245 ( .B1(n4333), .B2(n762), .C1(n4298), .C2(n219), .A(n854), 
        .ZN(U62_Z_66) );
  OAI221_X2 U247 ( .B1(n4333), .B2(n763), .C1(n4298), .C2(n220), .A(n856), 
        .ZN(U62_Z_65) );
  OAI221_X2 U249 ( .B1(n4333), .B2(n764), .C1(n4286), .C2(n221), .A(n858), 
        .ZN(U62_Z_64) );
  OAI221_X2 U255 ( .B1(n4302), .B2(n758), .C1(n4286), .C2(n263), .A(n866), 
        .ZN(U62_Z_6) );
  OAI221_X2 U267 ( .B1(n802), .B2(n759), .C1(n4286), .C2(n264), .A(n877), .ZN(
        U62_Z_5) );
  OAI221_X2 U271 ( .B1(n4302), .B2(n717), .C1(n4286), .C2(n222), .A(n880), 
        .ZN(U62_Z_47) );
  OAI221_X2 U273 ( .B1(n802), .B2(n718), .C1(n4286), .C2(n223), .A(n882), .ZN(
        U62_Z_46) );
  OAI221_X2 U275 ( .B1(n4302), .B2(n719), .C1(n4286), .C2(n224), .A(n884), 
        .ZN(U62_Z_45) );
  OAI221_X2 U277 ( .B1(n4302), .B2(n720), .C1(n4286), .C2(n225), .A(n886), 
        .ZN(U62_Z_44) );
  OAI221_X2 U279 ( .B1(n4302), .B2(n721), .C1(n4286), .C2(n226), .A(n888), 
        .ZN(U62_Z_43) );
  OAI221_X2 U281 ( .B1(n4302), .B2(n722), .C1(n4297), .C2(n227), .A(n890), 
        .ZN(U62_Z_42) );
  OAI221_X2 U283 ( .B1(n4302), .B2(n723), .C1(n4298), .C2(n228), .A(n892), 
        .ZN(U62_Z_41) );
  OAI221_X2 U285 ( .B1(n4302), .B2(n724), .C1(n4299), .C2(n229), .A(n894), 
        .ZN(U62_Z_40) );
  OAI221_X2 U287 ( .B1(n4302), .B2(n760), .C1(n4297), .C2(n265), .A(n896), 
        .ZN(U62_Z_4) );
  OAI221_X2 U289 ( .B1(n4302), .B2(n725), .C1(n4298), .C2(n230), .A(n897), 
        .ZN(U62_Z_39) );
  OAI221_X2 U291 ( .B1(n4302), .B2(n726), .C1(n4298), .C2(n231), .A(n899), 
        .ZN(U62_Z_38) );
  OAI221_X2 U293 ( .B1(n4302), .B2(n727), .C1(n4299), .C2(n232), .A(n901), 
        .ZN(U62_Z_37) );
  OAI221_X2 U295 ( .B1(n4302), .B2(n728), .C1(n4299), .C2(n233), .A(n903), 
        .ZN(U62_Z_36) );
  OAI221_X2 U305 ( .B1(n733), .B2(n802), .C1(n4286), .C2(n238), .A(n909), .ZN(
        U62_Z_31) );
  OAI221_X2 U307 ( .B1(n734), .B2(n802), .C1(n4286), .C2(n239), .A(n910), .ZN(
        U62_Z_30) );
  OAI221_X2 U309 ( .B1(n4302), .B2(n761), .C1(n4286), .C2(n266), .A(n911), 
        .ZN(U62_Z_3) );
  OAI221_X2 U311 ( .B1(n735), .B2(n802), .C1(n4286), .C2(n240), .A(n912), .ZN(
        U62_Z_29) );
  OAI221_X2 U313 ( .B1(n736), .B2(n802), .C1(n4286), .C2(n241), .A(n913), .ZN(
        U62_Z_28) );
  OAI221_X2 U315 ( .B1(n737), .B2(n802), .C1(n4286), .C2(n242), .A(n914), .ZN(
        U62_Z_27) );
  OAI221_X2 U317 ( .B1(n738), .B2(n802), .C1(n4297), .C2(n243), .A(n915), .ZN(
        U62_Z_26) );
  OAI221_X2 U325 ( .B1(n4302), .B2(n739), .C1(n4299), .C2(n244), .A(n922), 
        .ZN(U62_Z_25) );
  OAI221_X2 U337 ( .B1(n4302), .B2(n740), .C1(n4299), .C2(n245), .A(n933), 
        .ZN(U62_Z_24) );
  OAI221_X2 U349 ( .B1(n4302), .B2(n741), .C1(n4299), .C2(n246), .A(n946), 
        .ZN(U62_Z_23) );
  OAI221_X2 U361 ( .B1(n4302), .B2(n742), .C1(n4299), .C2(n247), .A(n957), 
        .ZN(U62_Z_22) );
  OAI221_X2 U373 ( .B1(n4302), .B2(n743), .C1(n4299), .C2(n248), .A(n968), 
        .ZN(U62_Z_21) );
  OAI221_X2 U385 ( .B1(n802), .B2(n744), .C1(n4299), .C2(n249), .A(n979), .ZN(
        U62_Z_20) );
  OAI221_X2 U387 ( .B1(n802), .B2(n762), .C1(n4299), .C2(n267), .A(n980), .ZN(
        U62_Z_2) );
  OAI22_X2 U397 ( .A1(n123), .A2(n990), .B1(n991), .B2(n992), .ZN(n989) );
  NOR2_X2 U398 ( .A1(n274), .A2(n993), .ZN(n991) );
  NOR3_X2 U399 ( .A1(n994), .A2(n995), .A3(n996), .ZN(n990) );
  OAI22_X2 U400 ( .A1(n998), .A2(n992), .B1(n123), .B2(n272), .ZN(n997) );
  NOR3_X2 U401 ( .A1(n270), .A2(n275), .A3(n271), .ZN(n998) );
  OAI221_X2 U404 ( .B1(n802), .B2(n745), .C1(n4299), .C2(n250), .A(n1002), 
        .ZN(U62_Z_19) );
  OAI221_X2 U416 ( .B1(n802), .B2(n746), .C1(n4297), .C2(n251), .A(n1013), 
        .ZN(U62_Z_18) );
  OAI221_X2 U430 ( .B1(n721), .B2(n1018), .C1(n4299), .C2(n130), .A(n1025), 
        .ZN(U62_Z_171) );
  OAI221_X2 U432 ( .B1(n722), .B2(n1018), .C1(n4299), .C2(n131), .A(n1026), 
        .ZN(U62_Z_170) );
  OAI221_X2 U434 ( .B1(n802), .B2(n747), .C1(n4299), .C2(n252), .A(n1027), 
        .ZN(U62_Z_17) );
  OAI221_X2 U436 ( .B1(n723), .B2(n1018), .C1(n4299), .C2(n132), .A(n1028), 
        .ZN(U62_Z_169) );
  OAI221_X2 U438 ( .B1(n724), .B2(n1018), .C1(n4299), .C2(n133), .A(n1029), 
        .ZN(U62_Z_168) );
  OAI221_X2 U440 ( .B1(n725), .B2(n1018), .C1(n4299), .C2(n134), .A(n1030), 
        .ZN(U62_Z_167) );
  OAI221_X2 U442 ( .B1(n726), .B2(n1018), .C1(n4299), .C2(n135), .A(n1031), 
        .ZN(U62_Z_166) );
  OAI221_X2 U444 ( .B1(n727), .B2(n1018), .C1(n4299), .C2(n136), .A(n1032), 
        .ZN(U62_Z_165) );
  OAI221_X2 U446 ( .B1(n728), .B2(n1018), .C1(n4299), .C2(n137), .A(n1033), 
        .ZN(U62_Z_164) );
  OAI221_X2 U448 ( .B1(n729), .B2(n1018), .C1(n4299), .C2(n138), .A(n1034), 
        .ZN(U62_Z_163) );
  OAI22_X2 U450 ( .A1(n407), .A2(n4317), .B1(n4320), .B2(n359), .ZN(n782) );
  OAI221_X2 U451 ( .B1(n730), .B2(n1018), .C1(n4299), .C2(n139), .A(n1035), 
        .ZN(U62_Z_162) );
  OAI22_X2 U453 ( .A1(n408), .A2(n4317), .B1(n4279), .B2(n360), .ZN(n785) );
  OAI221_X2 U454 ( .B1(n731), .B2(n1018), .C1(n4299), .C2(n140), .A(n1036), 
        .ZN(U62_Z_161) );
  OAI22_X2 U456 ( .A1(n409), .A2(n4317), .B1(n4279), .B2(n361), .ZN(n787) );
  OAI221_X2 U457 ( .B1(n732), .B2(n1018), .C1(n4286), .C2(n141), .A(n1037), 
        .ZN(U62_Z_160) );
  OAI22_X2 U459 ( .A1(n410), .A2(n4317), .B1(n4320), .B2(n362), .ZN(n789) );
  OAI221_X2 U460 ( .B1(n802), .B2(n748), .C1(n4286), .C2(n253), .A(n1038), 
        .ZN(U62_Z_16) );
  OAI221_X2 U462 ( .B1(n733), .B2(n4294), .C1(n4286), .C2(n142), .A(n1039), 
        .ZN(U62_Z_159) );
  OAI22_X2 U464 ( .A1(n411), .A2(n4317), .B1(n4320), .B2(n363), .ZN(n791) );
  OAI221_X2 U465 ( .B1(n734), .B2(n4294), .C1(n4286), .C2(n143), .A(n1040), 
        .ZN(U62_Z_158) );
  OAI22_X2 U467 ( .A1(n412), .A2(n4318), .B1(n4320), .B2(n364), .ZN(n793) );
  OAI221_X2 U468 ( .B1(n735), .B2(n4294), .C1(n4286), .C2(n144), .A(n1041), 
        .ZN(U62_Z_157) );
  OAI22_X2 U470 ( .A1(n413), .A2(n4317), .B1(n4279), .B2(n365), .ZN(n795) );
  OAI221_X2 U471 ( .B1(n736), .B2(n4294), .C1(n4286), .C2(n145), .A(n1042), 
        .ZN(U62_Z_156) );
  OAI22_X2 U473 ( .A1(n414), .A2(n4317), .B1(n4320), .B2(n366), .ZN(n797) );
  OAI221_X2 U474 ( .B1(n737), .B2(n4294), .C1(n4286), .C2(n146), .A(n1043), 
        .ZN(U62_Z_155) );
  OAI22_X2 U476 ( .A1(n415), .A2(n4317), .B1(n4320), .B2(n367), .ZN(n799) );
  OAI221_X2 U477 ( .B1(n738), .B2(n4294), .C1(n4286), .C2(n147), .A(n1044), 
        .ZN(U62_Z_154) );
  OAI22_X2 U479 ( .A1(n416), .A2(n4318), .B1(n4279), .B2(n368), .ZN(n801) );
  OAI221_X2 U480 ( .B1(n739), .B2(n4294), .C1(n4286), .C2(n148), .A(n1045), 
        .ZN(U62_Z_153) );
  OAI22_X2 U482 ( .A1(n417), .A2(n4317), .B1(n4320), .B2(n369), .ZN(n808) );
  OAI221_X2 U483 ( .B1(n740), .B2(n4294), .C1(n4286), .C2(n149), .A(n1046), 
        .ZN(U62_Z_152) );
  OAI22_X2 U485 ( .A1(n418), .A2(n4318), .B1(n4320), .B2(n370), .ZN(n810) );
  OAI221_X2 U486 ( .B1(n741), .B2(n4294), .C1(n4286), .C2(n150), .A(n1047), 
        .ZN(U62_Z_151) );
  OAI22_X2 U488 ( .A1(n419), .A2(n4318), .B1(n4320), .B2(n371), .ZN(n812) );
  OAI221_X2 U489 ( .B1(n742), .B2(n4294), .C1(n4286), .C2(n151), .A(n1048), 
        .ZN(U62_Z_150) );
  OAI22_X2 U491 ( .A1(n420), .A2(n4318), .B1(n4279), .B2(n372), .ZN(n814) );
  OAI221_X2 U492 ( .B1(n802), .B2(n749), .C1(n4299), .C2(n254), .A(n1049), 
        .ZN(U62_Z_15) );
  OAI221_X2 U494 ( .B1(n743), .B2(n4294), .C1(n4299), .C2(n152), .A(n1050), 
        .ZN(U62_Z_149) );
  OAI22_X2 U496 ( .A1(n421), .A2(n4318), .B1(n4320), .B2(n373), .ZN(n816) );
  OAI221_X2 U497 ( .B1(n744), .B2(n4294), .C1(n4297), .C2(n153), .A(n1051), 
        .ZN(U62_Z_148) );
  OAI22_X2 U499 ( .A1(n422), .A2(n4318), .B1(n4320), .B2(n374), .ZN(n818) );
  OAI221_X2 U500 ( .B1(n745), .B2(n4294), .C1(n4298), .C2(n154), .A(n1052), 
        .ZN(U62_Z_147) );
  OAI22_X2 U502 ( .A1(n423), .A2(n4318), .B1(n4320), .B2(n375), .ZN(n820) );
  OAI221_X2 U503 ( .B1(n746), .B2(n4294), .C1(n4286), .C2(n155), .A(n1053), 
        .ZN(U62_Z_146) );
  OAI22_X2 U505 ( .A1(n424), .A2(n4318), .B1(n4320), .B2(n376), .ZN(n822) );
  OAI221_X2 U506 ( .B1(n747), .B2(n4294), .C1(n4286), .C2(n156), .A(n1054), 
        .ZN(U62_Z_145) );
  OAI22_X2 U508 ( .A1(n425), .A2(n4318), .B1(n4320), .B2(n377), .ZN(n824) );
  OAI221_X2 U509 ( .B1(n748), .B2(n4294), .C1(n4286), .C2(n157), .A(n1055), 
        .ZN(U62_Z_144) );
  OAI22_X2 U511 ( .A1(n426), .A2(n4318), .B1(n4320), .B2(n378), .ZN(n826) );
  OAI221_X2 U512 ( .B1(n749), .B2(n4294), .C1(n4286), .C2(n158), .A(n1056), 
        .ZN(U62_Z_143) );
  OAI22_X2 U514 ( .A1(n427), .A2(n4318), .B1(n4320), .B2(n379), .ZN(n830) );
  OAI221_X2 U515 ( .B1(n750), .B2(n4294), .C1(n4286), .C2(n159), .A(n1057), 
        .ZN(U62_Z_142) );
  OAI221_X2 U517 ( .B1(n751), .B2(n4294), .C1(n4286), .C2(n160), .A(n1058), 
        .ZN(U62_Z_141) );
  OAI221_X2 U519 ( .B1(n752), .B2(n4294), .C1(n4286), .C2(n161), .A(n1059), 
        .ZN(U62_Z_140) );
  OAI221_X2 U521 ( .B1(n802), .B2(n750), .C1(n4286), .C2(n255), .A(n1060), 
        .ZN(U62_Z_14) );
  OAI22_X2 U523 ( .A1(n428), .A2(n4318), .B1(n4320), .B2(n380), .ZN(n832) );
  OAI221_X2 U524 ( .B1(n753), .B2(n4294), .C1(n4286), .C2(n162), .A(n1061), 
        .ZN(U62_Z_139) );
  OAI221_X2 U526 ( .B1(n754), .B2(n4294), .C1(n4286), .C2(n163), .A(n1062), 
        .ZN(U62_Z_138) );
  OAI221_X2 U528 ( .B1(n755), .B2(n4294), .C1(n4298), .C2(n164), .A(n1063), 
        .ZN(U62_Z_137) );
  OAI22_X2 U530 ( .A1(n433), .A2(n4318), .B1(n4320), .B2(n385), .ZN(n806) );
  OAI221_X2 U531 ( .B1(n756), .B2(n1018), .C1(n4299), .C2(n165), .A(n1064), 
        .ZN(U62_Z_136) );
  OAI22_X2 U533 ( .A1(n434), .A2(n4318), .B1(n4320), .B2(n386), .ZN(n828) );
  OAI221_X2 U534 ( .B1(n757), .B2(n4294), .C1(n4299), .C2(n166), .A(n1065), 
        .ZN(U62_Z_135) );
  OAI22_X2 U536 ( .A1(n435), .A2(n4318), .B1(n4320), .B2(n387), .ZN(n844) );
  OAI221_X2 U537 ( .B1(n758), .B2(n1018), .C1(n4298), .C2(n167), .A(n1066), 
        .ZN(U62_Z_134) );
  OAI22_X2 U539 ( .A1(n436), .A2(n4318), .B1(n4320), .B2(n388), .ZN(n846) );
  OAI221_X2 U540 ( .B1(n759), .B2(n4294), .C1(n4299), .C2(n168), .A(n1067), 
        .ZN(U62_Z_133) );
  OAI22_X2 U542 ( .A1(n437), .A2(n4318), .B1(n4279), .B2(n389), .ZN(n849) );
  OAI221_X2 U543 ( .B1(n760), .B2(n1018), .C1(n4298), .C2(n169), .A(n1068), 
        .ZN(U62_Z_132) );
  OAI22_X2 U545 ( .A1(n438), .A2(n4318), .B1(n4320), .B2(n390), .ZN(n851) );
  OAI221_X2 U546 ( .B1(n761), .B2(n4294), .C1(n4298), .C2(n170), .A(n1069), 
        .ZN(U62_Z_131) );
  OAI22_X2 U548 ( .A1(n439), .A2(n4318), .B1(n4320), .B2(n391), .ZN(n853) );
  OAI221_X2 U549 ( .B1(n762), .B2(n4294), .C1(n4298), .C2(n171), .A(n1070), 
        .ZN(U62_Z_130) );
  OAI22_X2 U551 ( .A1(n440), .A2(n4318), .B1(n4279), .B2(n392), .ZN(n855) );
  OAI221_X2 U552 ( .B1(n802), .B2(n751), .C1(n4298), .C2(n256), .A(n1071), 
        .ZN(U62_Z_13) );
  OAI22_X2 U554 ( .A1(n429), .A2(n4318), .B1(n4279), .B2(n381), .ZN(n834) );
  OAI221_X2 U555 ( .B1(n763), .B2(n1018), .C1(n4298), .C2(n172), .A(n1072), 
        .ZN(U62_Z_129) );
  OAI221_X2 U557 ( .B1(n764), .B2(n1018), .C1(n4298), .C2(n173), .A(n1073), 
        .ZN(U62_Z_128) );
  OAI22_X2 U559 ( .A1(n1075), .A2(n992), .B1(n123), .B2(n1076), .ZN(n1074) );
  NOR3_X2 U560 ( .A1(n994), .A2(n995), .A3(n999), .ZN(n1076) );
  NOR3_X2 U561 ( .A1(n274), .A2(n275), .A3(n270), .ZN(n1075) );
  NAND2_X2 U564 ( .A1(n1081), .A2(n1082), .ZN(n993) );
  NAND2_X2 U565 ( .A1(n271), .A2(n1083), .ZN(n1018) );
  OAI221_X2 U574 ( .B1(n4302), .B2(n752), .C1(n4298), .C2(n257), .A(n1092), 
        .ZN(U62_Z_12) );
  OAI22_X2 U576 ( .A1(n430), .A2(n4318), .B1(n4320), .B2(n382), .ZN(n836) );
  NOR3_X2 U587 ( .A1(n1105), .A2(n274), .A3(n1106), .ZN(n1102) );
  OAI221_X2 U588 ( .B1(n4333), .B2(n717), .C1(n4298), .C2(n174), .A(n1107), 
        .ZN(U62_Z_111) );
  OAI22_X2 U590 ( .A1(n395), .A2(n4317), .B1(n4320), .B2(n347), .ZN(n881) );
  OAI221_X2 U591 ( .B1(n4333), .B2(n718), .C1(n4299), .C2(n175), .A(n1108), 
        .ZN(U62_Z_110) );
  OAI22_X2 U593 ( .A1(n396), .A2(n4269), .B1(n4319), .B2(n348), .ZN(n883) );
  OAI221_X2 U594 ( .B1(n4302), .B2(n753), .C1(n4299), .C2(n258), .A(n1109), 
        .ZN(U62_Z_11) );
  OAI22_X2 U596 ( .A1(n431), .A2(n4317), .B1(n4320), .B2(n383), .ZN(n838) );
  OAI221_X2 U597 ( .B1(n4333), .B2(n719), .C1(n4299), .C2(n176), .A(n1110), 
        .ZN(U62_Z_109) );
  OAI22_X2 U599 ( .A1(n397), .A2(n4317), .B1(n4320), .B2(n349), .ZN(n885) );
  OAI221_X2 U600 ( .B1(n4333), .B2(n720), .C1(n4299), .C2(n177), .A(n1111), 
        .ZN(U62_Z_108) );
  OAI22_X2 U602 ( .A1(n398), .A2(n4269), .B1(n4320), .B2(n350), .ZN(n887) );
  OAI221_X2 U603 ( .B1(n4333), .B2(n721), .C1(n4299), .C2(n178), .A(n1112), 
        .ZN(U62_Z_107) );
  OAI22_X2 U605 ( .A1(n399), .A2(n4317), .B1(n4320), .B2(n351), .ZN(n889) );
  OAI221_X2 U606 ( .B1(n4333), .B2(n722), .C1(n4299), .C2(n179), .A(n1113), 
        .ZN(U62_Z_106) );
  OAI22_X2 U608 ( .A1(n400), .A2(n4317), .B1(n4320), .B2(n352), .ZN(n891) );
  OAI221_X2 U609 ( .B1(n4333), .B2(n723), .C1(n4299), .C2(n180), .A(n1114), 
        .ZN(U62_Z_105) );
  OAI22_X2 U611 ( .A1(n401), .A2(n4269), .B1(n4320), .B2(n353), .ZN(n893) );
  OAI221_X2 U612 ( .B1(n4333), .B2(n724), .C1(n4299), .C2(n181), .A(n1115), 
        .ZN(U62_Z_104) );
  OAI22_X2 U614 ( .A1(n402), .A2(n4317), .B1(n4320), .B2(n354), .ZN(n895) );
  OAI221_X2 U615 ( .B1(n4333), .B2(n725), .C1(n4299), .C2(n182), .A(n1116), 
        .ZN(U62_Z_103) );
  OAI22_X2 U617 ( .A1(n403), .A2(n4317), .B1(n4320), .B2(n355), .ZN(n898) );
  OAI221_X2 U618 ( .B1(n4333), .B2(n726), .C1(n4298), .C2(n183), .A(n1117), 
        .ZN(U62_Z_102) );
  OAI22_X2 U620 ( .A1(n404), .A2(n4269), .B1(n4320), .B2(n356), .ZN(n900) );
  OAI221_X2 U621 ( .B1(n4333), .B2(n727), .C1(n4298), .C2(n184), .A(n1118), 
        .ZN(U62_Z_101) );
  OAI22_X2 U623 ( .A1(n405), .A2(n4317), .B1(n4320), .B2(n357), .ZN(n902) );
  OAI221_X2 U624 ( .B1(n4333), .B2(n728), .C1(n4299), .C2(n185), .A(n1119), 
        .ZN(U62_Z_100) );
  NOR2_X2 U626 ( .A1(n1079), .A2(n1120), .ZN(n783) );
  NAND3_X2 U628 ( .A1(n1121), .A2(n1081), .A3(n1077), .ZN(n1105) );
  OAI22_X2 U629 ( .A1(n406), .A2(n4317), .B1(n4320), .B2(n358), .ZN(n904) );
  OAI221_X2 U633 ( .B1(n4302), .B2(n754), .C1(n4298), .C2(n259), .A(n1124), 
        .ZN(U62_Z_10) );
  OAI22_X2 U635 ( .A1(n432), .A2(n4269), .B1(n4320), .B2(n384), .ZN(n840) );
  OAI221_X2 U636 ( .B1(n4302), .B2(n763), .C1(n4299), .C2(n268), .A(n1125), 
        .ZN(U62_Z_1) );
  OAI22_X2 U638 ( .A1(n441), .A2(n4317), .B1(n4320), .B2(n393), .ZN(n857) );
  OAI221_X2 U639 ( .B1(n802), .B2(n764), .C1(n4299), .C2(n269), .A(n1126), 
        .ZN(U62_Z_0) );
  OAI22_X2 U641 ( .A1(n442), .A2(n4317), .B1(n4320), .B2(n394), .ZN(n859) );
  NOR4_X2 U642 ( .A1(n273), .A2(n277), .A3(n276), .A4(n1128), .ZN(n995) );
  OAI22_X2 U643 ( .A1(n123), .A2(n1130), .B1(n1131), .B2(n992), .ZN(n1129) );
  NOR2_X2 U644 ( .A1(n271), .A2(n1106), .ZN(n1131) );
  NAND2_X2 U645 ( .A1(n1082), .A2(n1078), .ZN(n1106) );
  NAND3_X2 U646 ( .A1(n1132), .A2(n1133), .A3(n1134), .ZN(n1078) );
  NAND3_X2 U648 ( .A1(n1137), .A2(n1138), .A3(n1139), .ZN(n1082) );
  NAND2_X2 U650 ( .A1(n1132), .A2(n1141), .ZN(n1121) );
  NOR3_X2 U652 ( .A1(n994), .A2(n996), .A3(n999), .ZN(n1130) );
  NOR4_X2 U653 ( .A1(n273), .A2(n277), .A3(n278), .A4(n1142), .ZN(n999) );
  NOR4_X2 U654 ( .A1(n273), .A2(n278), .A3(n276), .A4(n1140), .ZN(n996) );
  NOR4_X2 U655 ( .A1(n277), .A2(n278), .A3(n276), .A4(n1136), .ZN(n994) );
  NAND2_X2 U656 ( .A1(n1083), .A2(n1144), .ZN(n802) );
  NAND3_X2 U657 ( .A1(n1077), .A2(n1081), .A3(n1123), .ZN(n1144) );
  NAND2_X2 U658 ( .A1(n1137), .A2(n1145), .ZN(n1123) );
  NAND3_X2 U660 ( .A1(n1141), .A2(n1143), .A3(n1146), .ZN(n1081) );
  NAND3_X2 U663 ( .A1(n1145), .A2(n1135), .A3(n1147), .ZN(n1077) );
  OAI221_X2 U670 ( .B1(n1148), .B2(n4297), .C1(n4290), .C2(n1150), .A(n5), 
        .ZN(U61_Z_9) );
  OAI221_X2 U671 ( .B1(n1151), .B2(n4297), .C1(n4290), .C2(n1152), .A(n5), 
        .ZN(U61_Z_8) );
  OAI221_X2 U672 ( .B1(n1153), .B2(n4297), .C1(n4290), .C2(n1154), .A(n5), 
        .ZN(U61_Z_7) );
  OAI221_X2 U673 ( .B1(n1155), .B2(n4297), .C1(n4290), .C2(n1156), .A(n5), 
        .ZN(U61_Z_6) );
  OAI221_X2 U674 ( .B1(n1157), .B2(n4297), .C1(n4290), .C2(n1158), .A(n5), 
        .ZN(U61_Z_5) );
  OAI221_X2 U675 ( .B1(n1159), .B2(n4298), .C1(n4290), .C2(n1160), .A(n5), 
        .ZN(U61_Z_4) );
  OAI221_X2 U676 ( .B1(n1161), .B2(n4297), .C1(n4290), .C2(n1162), .A(n5), 
        .ZN(U61_Z_3) );
  OAI221_X2 U677 ( .B1(n1163), .B2(n4297), .C1(n4290), .C2(n1164), .A(n5), 
        .ZN(U61_Z_2) );
  OAI221_X2 U678 ( .B1(n1165), .B2(n4297), .C1(n4290), .C2(n1166), .A(n5), 
        .ZN(U61_Z_10) );
  OAI221_X2 U679 ( .B1(n1167), .B2(n4297), .C1(n4290), .C2(n1168), .A(n5), 
        .ZN(U61_Z_1) );
  OAI221_X2 U680 ( .B1(n1169), .B2(n4297), .C1(n4290), .C2(n1170), .A(n5), 
        .ZN(U61_Z_0) );
  NAND3_X2 U693 ( .A1(n778), .A2(n772), .A3(n992), .ZN(n1182) );
  NOR2_X2 U694 ( .A1(n774), .A2(n4318), .ZN(U58_Z_0) );
  NOR2_X2 U695 ( .A1(n4296), .A2(n1083), .ZN(n774) );
  NOR2_X2 U696 ( .A1(n1079), .A2(n992), .ZN(n1083) );
  OAI22_X2 U697 ( .A1(n729), .A2(n4325), .B1(n4278), .B2(n585), .ZN(U57_Z_99)
         );
  OAI22_X2 U698 ( .A1(n730), .A2(n4325), .B1(n4278), .B2(n586), .ZN(U57_Z_98)
         );
  OAI22_X2 U699 ( .A1(n731), .A2(n4325), .B1(n4278), .B2(n587), .ZN(U57_Z_97)
         );
  OAI22_X2 U700 ( .A1(n732), .A2(n4325), .B1(n4278), .B2(n588), .ZN(U57_Z_96)
         );
  OAI22_X2 U701 ( .A1(n733), .A2(n4325), .B1(n4278), .B2(n589), .ZN(U57_Z_95)
         );
  OAI22_X2 U702 ( .A1(n734), .A2(n4325), .B1(n4278), .B2(n590), .ZN(U57_Z_94)
         );
  OAI22_X2 U703 ( .A1(n735), .A2(n4325), .B1(n4278), .B2(n591), .ZN(U57_Z_93)
         );
  OAI22_X2 U704 ( .A1(n736), .A2(n4325), .B1(n4278), .B2(n592), .ZN(U57_Z_92)
         );
  OAI22_X2 U705 ( .A1(n737), .A2(n4325), .B1(n4278), .B2(n593), .ZN(U57_Z_91)
         );
  OAI22_X2 U706 ( .A1(n738), .A2(n4325), .B1(n4278), .B2(n594), .ZN(U57_Z_90)
         );
  OAI22_X2 U707 ( .A1(n755), .A2(n4327), .B1(n4277), .B2(n659), .ZN(U57_Z_9)
         );
  OAI22_X2 U708 ( .A1(n739), .A2(n4325), .B1(n4278), .B2(n595), .ZN(U57_Z_89)
         );
  OAI22_X2 U709 ( .A1(n740), .A2(n4325), .B1(n4278), .B2(n596), .ZN(U57_Z_88)
         );
  OAI22_X2 U710 ( .A1(n741), .A2(n4325), .B1(n4278), .B2(n597), .ZN(U57_Z_87)
         );
  OAI22_X2 U711 ( .A1(n742), .A2(n4325), .B1(n4278), .B2(n598), .ZN(U57_Z_86)
         );
  OAI22_X2 U712 ( .A1(n743), .A2(n4325), .B1(n4278), .B2(n599), .ZN(U57_Z_85)
         );
  OAI22_X2 U713 ( .A1(n744), .A2(n4325), .B1(n4278), .B2(n600), .ZN(U57_Z_84)
         );
  OAI22_X2 U714 ( .A1(n745), .A2(n4325), .B1(n4278), .B2(n601), .ZN(U57_Z_83)
         );
  OAI22_X2 U715 ( .A1(n746), .A2(n4325), .B1(n4278), .B2(n602), .ZN(U57_Z_82)
         );
  OAI22_X2 U716 ( .A1(n747), .A2(n4325), .B1(n4278), .B2(n603), .ZN(U57_Z_81)
         );
  OAI22_X2 U717 ( .A1(n748), .A2(n4325), .B1(n4278), .B2(n604), .ZN(U57_Z_80)
         );
  OAI22_X2 U718 ( .A1(n756), .A2(n4327), .B1(n4277), .B2(n660), .ZN(U57_Z_8)
         );
  OAI22_X2 U719 ( .A1(n749), .A2(n4325), .B1(n4278), .B2(n605), .ZN(U57_Z_79)
         );
  OAI22_X2 U720 ( .A1(n750), .A2(n4325), .B1(n4278), .B2(n606), .ZN(U57_Z_78)
         );
  OAI22_X2 U721 ( .A1(n751), .A2(n4325), .B1(n4278), .B2(n607), .ZN(U57_Z_77)
         );
  OAI22_X2 U722 ( .A1(n752), .A2(n4325), .B1(n4278), .B2(n608), .ZN(U57_Z_76)
         );
  OAI22_X2 U723 ( .A1(n753), .A2(n4325), .B1(n4278), .B2(n609), .ZN(U57_Z_75)
         );
  OAI22_X2 U724 ( .A1(n754), .A2(n4325), .B1(n4278), .B2(n610), .ZN(U57_Z_74)
         );
  OAI22_X2 U725 ( .A1(n755), .A2(n4325), .B1(n4278), .B2(n611), .ZN(U57_Z_73)
         );
  OAI22_X2 U726 ( .A1(n756), .A2(n4325), .B1(n4278), .B2(n612), .ZN(U57_Z_72)
         );
  OAI22_X2 U727 ( .A1(n757), .A2(n4325), .B1(n4278), .B2(n613), .ZN(U57_Z_71)
         );
  OAI22_X2 U728 ( .A1(n758), .A2(n4325), .B1(n4278), .B2(n614), .ZN(U57_Z_70)
         );
  OAI22_X2 U729 ( .A1(n757), .A2(n4327), .B1(n4277), .B2(n661), .ZN(U57_Z_7)
         );
  OAI22_X2 U730 ( .A1(n759), .A2(n4325), .B1(n4278), .B2(n615), .ZN(U57_Z_69)
         );
  OAI22_X2 U731 ( .A1(n760), .A2(n4325), .B1(n4278), .B2(n616), .ZN(U57_Z_68)
         );
  OAI22_X2 U732 ( .A1(n761), .A2(n4325), .B1(n4278), .B2(n617), .ZN(U57_Z_67)
         );
  OAI22_X2 U733 ( .A1(n762), .A2(n4325), .B1(n4278), .B2(n618), .ZN(U57_Z_66)
         );
  OAI22_X2 U734 ( .A1(n763), .A2(n4325), .B1(n4278), .B2(n619), .ZN(U57_Z_65)
         );
  OAI22_X2 U735 ( .A1(n764), .A2(n4325), .B1(n4278), .B2(n620), .ZN(U57_Z_64)
         );
  OAI22_X2 U736 ( .A1(n758), .A2(n4327), .B1(n4277), .B2(n662), .ZN(U57_Z_6)
         );
  OAI22_X2 U737 ( .A1(n759), .A2(n4327), .B1(n4277), .B2(n663), .ZN(U57_Z_5)
         );
  OAI22_X2 U738 ( .A1(n717), .A2(n4327), .B1(n4277), .B2(n621), .ZN(U57_Z_47)
         );
  OAI22_X2 U739 ( .A1(n718), .A2(n4327), .B1(n4277), .B2(n622), .ZN(U57_Z_46)
         );
  OAI22_X2 U740 ( .A1(n719), .A2(n4327), .B1(n4277), .B2(n623), .ZN(U57_Z_45)
         );
  OAI22_X2 U741 ( .A1(n720), .A2(n4327), .B1(n4277), .B2(n624), .ZN(U57_Z_44)
         );
  OAI22_X2 U742 ( .A1(n721), .A2(n4327), .B1(n4277), .B2(n625), .ZN(U57_Z_43)
         );
  OAI22_X2 U743 ( .A1(n722), .A2(n4327), .B1(n4277), .B2(n626), .ZN(U57_Z_42)
         );
  OAI22_X2 U744 ( .A1(n723), .A2(n4327), .B1(n4277), .B2(n627), .ZN(U57_Z_41)
         );
  OAI22_X2 U745 ( .A1(n724), .A2(n4327), .B1(n4277), .B2(n628), .ZN(U57_Z_40)
         );
  OAI22_X2 U746 ( .A1(n760), .A2(n4327), .B1(n4277), .B2(n664), .ZN(U57_Z_4)
         );
  OAI22_X2 U747 ( .A1(n725), .A2(n4327), .B1(n4277), .B2(n629), .ZN(U57_Z_39)
         );
  OAI22_X2 U748 ( .A1(n726), .A2(n4327), .B1(n4277), .B2(n630), .ZN(U57_Z_38)
         );
  OAI22_X2 U749 ( .A1(n727), .A2(n4327), .B1(n4277), .B2(n631), .ZN(U57_Z_37)
         );
  OAI22_X2 U750 ( .A1(n728), .A2(n4327), .B1(n4277), .B2(n632), .ZN(U57_Z_36)
         );
  OAI22_X2 U751 ( .A1(n729), .A2(n4327), .B1(n4277), .B2(n633), .ZN(U57_Z_35)
         );
  OAI22_X2 U752 ( .A1(n730), .A2(n4327), .B1(n4277), .B2(n634), .ZN(U57_Z_34)
         );
  OAI22_X2 U753 ( .A1(n731), .A2(n4327), .B1(n4277), .B2(n635), .ZN(U57_Z_33)
         );
  OAI22_X2 U754 ( .A1(n732), .A2(n4327), .B1(n4277), .B2(n636), .ZN(U57_Z_32)
         );
  OAI22_X2 U755 ( .A1(n733), .A2(n4327), .B1(n4277), .B2(n637), .ZN(U57_Z_31)
         );
  OAI22_X2 U756 ( .A1(n734), .A2(n4327), .B1(n4277), .B2(n638), .ZN(U57_Z_30)
         );
  OAI22_X2 U757 ( .A1(n761), .A2(n4327), .B1(n4277), .B2(n665), .ZN(U57_Z_3)
         );
  OAI22_X2 U758 ( .A1(n735), .A2(n4327), .B1(n4277), .B2(n639), .ZN(U57_Z_29)
         );
  OAI22_X2 U759 ( .A1(n736), .A2(n4327), .B1(n4277), .B2(n640), .ZN(U57_Z_28)
         );
  OAI22_X2 U760 ( .A1(n737), .A2(n4327), .B1(n4277), .B2(n641), .ZN(U57_Z_27)
         );
  OAI22_X2 U761 ( .A1(n738), .A2(n4327), .B1(n4277), .B2(n642), .ZN(U57_Z_26)
         );
  OAI22_X2 U762 ( .A1(n739), .A2(n4327), .B1(n4277), .B2(n643), .ZN(U57_Z_25)
         );
  OAI22_X2 U763 ( .A1(n740), .A2(n4327), .B1(n4277), .B2(n644), .ZN(U57_Z_24)
         );
  OAI22_X2 U764 ( .A1(n717), .A2(n4329), .B1(n4273), .B2(n477), .ZN(U57_Z_239)
         );
  OAI22_X2 U765 ( .A1(n718), .A2(n4329), .B1(n4273), .B2(n478), .ZN(U57_Z_238)
         );
  OAI22_X2 U766 ( .A1(n719), .A2(n4329), .B1(n4273), .B2(n479), .ZN(U57_Z_237)
         );
  OAI22_X2 U767 ( .A1(n720), .A2(n4329), .B1(n4273), .B2(n480), .ZN(U57_Z_236)
         );
  OAI22_X2 U768 ( .A1(n721), .A2(n4329), .B1(n4273), .B2(n481), .ZN(U57_Z_235)
         );
  OAI22_X2 U769 ( .A1(n722), .A2(n4329), .B1(n4273), .B2(n482), .ZN(U57_Z_234)
         );
  OAI22_X2 U770 ( .A1(n723), .A2(n4329), .B1(n4273), .B2(n483), .ZN(U57_Z_233)
         );
  OAI22_X2 U771 ( .A1(n724), .A2(n4329), .B1(n4273), .B2(n484), .ZN(U57_Z_232)
         );
  OAI22_X2 U772 ( .A1(n725), .A2(n4329), .B1(n4273), .B2(n485), .ZN(U57_Z_231)
         );
  OAI22_X2 U773 ( .A1(n726), .A2(n4329), .B1(n4273), .B2(n486), .ZN(U57_Z_230)
         );
  OAI22_X2 U774 ( .A1(n741), .A2(n4327), .B1(n4277), .B2(n645), .ZN(U57_Z_23)
         );
  OAI22_X2 U775 ( .A1(n727), .A2(n4329), .B1(n4273), .B2(n487), .ZN(U57_Z_229)
         );
  OAI22_X2 U776 ( .A1(n728), .A2(n4329), .B1(n4273), .B2(n488), .ZN(U57_Z_228)
         );
  OAI22_X2 U777 ( .A1(n729), .A2(n4329), .B1(n4273), .B2(n489), .ZN(U57_Z_227)
         );
  OAI22_X2 U778 ( .A1(n730), .A2(n4329), .B1(n4273), .B2(n490), .ZN(U57_Z_226)
         );
  OAI22_X2 U779 ( .A1(n731), .A2(n4329), .B1(n4273), .B2(n491), .ZN(U57_Z_225)
         );
  OAI22_X2 U780 ( .A1(n732), .A2(n4329), .B1(n4273), .B2(n492), .ZN(U57_Z_224)
         );
  OAI22_X2 U781 ( .A1(n733), .A2(n4329), .B1(n4273), .B2(n493), .ZN(U57_Z_223)
         );
  OAI22_X2 U782 ( .A1(n734), .A2(n4329), .B1(n4273), .B2(n494), .ZN(U57_Z_222)
         );
  OAI22_X2 U783 ( .A1(n735), .A2(n4329), .B1(n4273), .B2(n495), .ZN(U57_Z_221)
         );
  OAI22_X2 U784 ( .A1(n736), .A2(n4329), .B1(n4273), .B2(n496), .ZN(U57_Z_220)
         );
  OAI22_X2 U785 ( .A1(n742), .A2(n4327), .B1(n4277), .B2(n646), .ZN(U57_Z_22)
         );
  OAI22_X2 U786 ( .A1(n737), .A2(n4329), .B1(n4273), .B2(n497), .ZN(U57_Z_219)
         );
  OAI22_X2 U787 ( .A1(n738), .A2(n4329), .B1(n4273), .B2(n498), .ZN(U57_Z_218)
         );
  OAI22_X2 U788 ( .A1(n739), .A2(n4329), .B1(n4273), .B2(n499), .ZN(U57_Z_217)
         );
  OAI22_X2 U789 ( .A1(n740), .A2(n4329), .B1(n4273), .B2(n500), .ZN(U57_Z_216)
         );
  OAI22_X2 U790 ( .A1(n741), .A2(n4329), .B1(n4273), .B2(n501), .ZN(U57_Z_215)
         );
  OAI22_X2 U791 ( .A1(n742), .A2(n4329), .B1(n4273), .B2(n502), .ZN(U57_Z_214)
         );
  OAI22_X2 U792 ( .A1(n743), .A2(n4329), .B1(n4273), .B2(n503), .ZN(U57_Z_213)
         );
  OAI22_X2 U793 ( .A1(n744), .A2(n4329), .B1(n4273), .B2(n504), .ZN(U57_Z_212)
         );
  OAI22_X2 U794 ( .A1(n745), .A2(n4329), .B1(n4273), .B2(n505), .ZN(U57_Z_211)
         );
  OAI22_X2 U795 ( .A1(n746), .A2(n4329), .B1(n4273), .B2(n506), .ZN(U57_Z_210)
         );
  OAI22_X2 U796 ( .A1(n743), .A2(n4327), .B1(n4277), .B2(n647), .ZN(U57_Z_21)
         );
  OAI22_X2 U797 ( .A1(n747), .A2(n4329), .B1(n4273), .B2(n507), .ZN(U57_Z_209)
         );
  OAI22_X2 U798 ( .A1(n748), .A2(n4329), .B1(n4273), .B2(n508), .ZN(U57_Z_208)
         );
  OAI22_X2 U799 ( .A1(n749), .A2(n4329), .B1(n4273), .B2(n509), .ZN(U57_Z_207)
         );
  OAI22_X2 U800 ( .A1(n750), .A2(n4329), .B1(n4273), .B2(n510), .ZN(U57_Z_206)
         );
  OAI22_X2 U801 ( .A1(n751), .A2(n4329), .B1(n4273), .B2(n511), .ZN(U57_Z_205)
         );
  OAI22_X2 U802 ( .A1(n752), .A2(n4329), .B1(n4273), .B2(n512), .ZN(U57_Z_204)
         );
  OAI22_X2 U803 ( .A1(n753), .A2(n4329), .B1(n4273), .B2(n513), .ZN(U57_Z_203)
         );
  OAI22_X2 U804 ( .A1(n754), .A2(n4329), .B1(n4273), .B2(n514), .ZN(U57_Z_202)
         );
  OAI22_X2 U805 ( .A1(n755), .A2(n4329), .B1(n4273), .B2(n515), .ZN(U57_Z_201)
         );
  OAI22_X2 U806 ( .A1(n756), .A2(n4329), .B1(n4273), .B2(n516), .ZN(U57_Z_200)
         );
  OAI22_X2 U807 ( .A1(n744), .A2(n4327), .B1(n4277), .B2(n648), .ZN(U57_Z_20)
         );
  OAI22_X2 U808 ( .A1(n762), .A2(n4327), .B1(n4277), .B2(n666), .ZN(U57_Z_2)
         );
  OAI22_X2 U809 ( .A1(n757), .A2(n4329), .B1(n4273), .B2(n517), .ZN(U57_Z_199)
         );
  OAI22_X2 U810 ( .A1(n758), .A2(n4329), .B1(n4273), .B2(n518), .ZN(U57_Z_198)
         );
  OAI22_X2 U811 ( .A1(n759), .A2(n4329), .B1(n4273), .B2(n519), .ZN(U57_Z_197)
         );
  OAI22_X2 U812 ( .A1(n760), .A2(n4329), .B1(n4273), .B2(n520), .ZN(U57_Z_196)
         );
  OAI22_X2 U813 ( .A1(n761), .A2(n4329), .B1(n4273), .B2(n521), .ZN(U57_Z_195)
         );
  OAI22_X2 U814 ( .A1(n762), .A2(n4329), .B1(n4273), .B2(n522), .ZN(U57_Z_194)
         );
  OAI22_X2 U815 ( .A1(n763), .A2(n4329), .B1(n4273), .B2(n523), .ZN(U57_Z_193)
         );
  OAI22_X2 U816 ( .A1(n764), .A2(n4329), .B1(n4273), .B2(n524), .ZN(U57_Z_192)
         );
  NAND3_X2 U818 ( .A1(n279), .A2(n1191), .A3(n280), .ZN(n1190) );
  OAI22_X2 U820 ( .A1(n745), .A2(n4327), .B1(n4277), .B2(n649), .ZN(U57_Z_19)
         );
  OAI22_X2 U821 ( .A1(n746), .A2(n4327), .B1(n4277), .B2(n650), .ZN(U57_Z_18)
         );
  OAI22_X2 U822 ( .A1(n717), .A2(n4331), .B1(n4272), .B2(n525), .ZN(U57_Z_175)
         );
  OAI22_X2 U823 ( .A1(n718), .A2(n4331), .B1(n4272), .B2(n526), .ZN(U57_Z_174)
         );
  OAI22_X2 U824 ( .A1(n719), .A2(n4331), .B1(n4272), .B2(n527), .ZN(U57_Z_173)
         );
  OAI22_X2 U825 ( .A1(n720), .A2(n4331), .B1(n4272), .B2(n528), .ZN(U57_Z_172)
         );
  OAI22_X2 U826 ( .A1(n721), .A2(n4331), .B1(n4272), .B2(n529), .ZN(U57_Z_171)
         );
  OAI22_X2 U827 ( .A1(n722), .A2(n4331), .B1(n4272), .B2(n530), .ZN(U57_Z_170)
         );
  OAI22_X2 U828 ( .A1(n747), .A2(n4327), .B1(n4277), .B2(n651), .ZN(U57_Z_17)
         );
  OAI22_X2 U829 ( .A1(n723), .A2(n4331), .B1(n4272), .B2(n531), .ZN(U57_Z_169)
         );
  OAI22_X2 U830 ( .A1(n724), .A2(n4331), .B1(n4272), .B2(n532), .ZN(U57_Z_168)
         );
  OAI22_X2 U831 ( .A1(n725), .A2(n4331), .B1(n4272), .B2(n533), .ZN(U57_Z_167)
         );
  OAI22_X2 U832 ( .A1(n726), .A2(n4331), .B1(n4272), .B2(n534), .ZN(U57_Z_166)
         );
  OAI22_X2 U833 ( .A1(n727), .A2(n4331), .B1(n4272), .B2(n535), .ZN(U57_Z_165)
         );
  OAI22_X2 U834 ( .A1(n728), .A2(n4331), .B1(n4272), .B2(n536), .ZN(U57_Z_164)
         );
  OAI22_X2 U835 ( .A1(n729), .A2(n4331), .B1(n4272), .B2(n537), .ZN(U57_Z_163)
         );
  OAI22_X2 U836 ( .A1(n730), .A2(n4331), .B1(n4272), .B2(n538), .ZN(U57_Z_162)
         );
  OAI22_X2 U837 ( .A1(n731), .A2(n4331), .B1(n4272), .B2(n539), .ZN(U57_Z_161)
         );
  OAI22_X2 U838 ( .A1(n732), .A2(n4331), .B1(n4272), .B2(n540), .ZN(U57_Z_160)
         );
  OAI22_X2 U839 ( .A1(n748), .A2(n4327), .B1(n4277), .B2(n652), .ZN(U57_Z_16)
         );
  OAI22_X2 U840 ( .A1(n733), .A2(n4331), .B1(n4272), .B2(n541), .ZN(U57_Z_159)
         );
  OAI22_X2 U841 ( .A1(n734), .A2(n4331), .B1(n4272), .B2(n542), .ZN(U57_Z_158)
         );
  OAI22_X2 U842 ( .A1(n735), .A2(n4331), .B1(n4272), .B2(n543), .ZN(U57_Z_157)
         );
  OAI22_X2 U843 ( .A1(n736), .A2(n4331), .B1(n4272), .B2(n544), .ZN(U57_Z_156)
         );
  OAI22_X2 U844 ( .A1(n737), .A2(n4331), .B1(n4272), .B2(n545), .ZN(U57_Z_155)
         );
  OAI22_X2 U845 ( .A1(n738), .A2(n4331), .B1(n4272), .B2(n546), .ZN(U57_Z_154)
         );
  OAI22_X2 U846 ( .A1(n739), .A2(n4331), .B1(n4272), .B2(n547), .ZN(U57_Z_153)
         );
  OAI22_X2 U847 ( .A1(n740), .A2(n4331), .B1(n4272), .B2(n548), .ZN(U57_Z_152)
         );
  OAI22_X2 U848 ( .A1(n741), .A2(n4331), .B1(n4272), .B2(n549), .ZN(U57_Z_151)
         );
  OAI22_X2 U849 ( .A1(n742), .A2(n4331), .B1(n4272), .B2(n550), .ZN(U57_Z_150)
         );
  OAI22_X2 U850 ( .A1(n749), .A2(n4327), .B1(n4277), .B2(n653), .ZN(U57_Z_15)
         );
  OAI22_X2 U851 ( .A1(n743), .A2(n4331), .B1(n4272), .B2(n551), .ZN(U57_Z_149)
         );
  OAI22_X2 U852 ( .A1(n744), .A2(n4331), .B1(n4272), .B2(n552), .ZN(U57_Z_148)
         );
  OAI22_X2 U853 ( .A1(n745), .A2(n4331), .B1(n4272), .B2(n553), .ZN(U57_Z_147)
         );
  OAI22_X2 U854 ( .A1(n746), .A2(n4331), .B1(n4272), .B2(n554), .ZN(U57_Z_146)
         );
  OAI22_X2 U855 ( .A1(n747), .A2(n4331), .B1(n4272), .B2(n555), .ZN(U57_Z_145)
         );
  OAI22_X2 U856 ( .A1(n748), .A2(n4331), .B1(n4272), .B2(n556), .ZN(U57_Z_144)
         );
  OAI22_X2 U857 ( .A1(n749), .A2(n4331), .B1(n4272), .B2(n557), .ZN(U57_Z_143)
         );
  OAI22_X2 U858 ( .A1(n750), .A2(n4331), .B1(n4272), .B2(n558), .ZN(U57_Z_142)
         );
  OAI22_X2 U859 ( .A1(n751), .A2(n4331), .B1(n4272), .B2(n559), .ZN(U57_Z_141)
         );
  OAI22_X2 U860 ( .A1(n752), .A2(n4331), .B1(n4272), .B2(n560), .ZN(U57_Z_140)
         );
  OAI22_X2 U861 ( .A1(n750), .A2(n4327), .B1(n4277), .B2(n654), .ZN(U57_Z_14)
         );
  OAI22_X2 U862 ( .A1(n753), .A2(n4331), .B1(n4272), .B2(n561), .ZN(U57_Z_139)
         );
  OAI22_X2 U863 ( .A1(n754), .A2(n4331), .B1(n4272), .B2(n562), .ZN(U57_Z_138)
         );
  OAI22_X2 U864 ( .A1(n755), .A2(n4331), .B1(n4272), .B2(n563), .ZN(U57_Z_137)
         );
  OAI22_X2 U865 ( .A1(n756), .A2(n4331), .B1(n4272), .B2(n564), .ZN(U57_Z_136)
         );
  OAI22_X2 U866 ( .A1(n757), .A2(n4331), .B1(n4272), .B2(n565), .ZN(U57_Z_135)
         );
  OAI22_X2 U867 ( .A1(n758), .A2(n4331), .B1(n4272), .B2(n566), .ZN(U57_Z_134)
         );
  OAI22_X2 U868 ( .A1(n759), .A2(n4331), .B1(n4272), .B2(n567), .ZN(U57_Z_133)
         );
  OAI22_X2 U869 ( .A1(n760), .A2(n4331), .B1(n4272), .B2(n568), .ZN(U57_Z_132)
         );
  OAI22_X2 U870 ( .A1(n761), .A2(n4331), .B1(n4272), .B2(n569), .ZN(U57_Z_131)
         );
  OAI22_X2 U871 ( .A1(n762), .A2(n4331), .B1(n4272), .B2(n570), .ZN(U57_Z_130)
         );
  OAI22_X2 U872 ( .A1(n751), .A2(n4327), .B1(n4277), .B2(n655), .ZN(U57_Z_13)
         );
  OAI22_X2 U873 ( .A1(n763), .A2(n4331), .B1(n4272), .B2(n571), .ZN(U57_Z_129)
         );
  OAI22_X2 U874 ( .A1(n764), .A2(n4331), .B1(n4272), .B2(n572), .ZN(U57_Z_128)
         );
  NAND3_X2 U876 ( .A1(n279), .A2(n1191), .A3(n281), .ZN(n1195) );
  OAI22_X2 U878 ( .A1(n752), .A2(n4327), .B1(n4277), .B2(n656), .ZN(U57_Z_12)
         );
  OAI22_X2 U880 ( .A1(n717), .A2(n4325), .B1(n4278), .B2(n573), .ZN(U57_Z_111)
         );
  OAI22_X2 U881 ( .A1(n718), .A2(n4325), .B1(n4278), .B2(n574), .ZN(U57_Z_110)
         );
  OAI22_X2 U882 ( .A1(n753), .A2(n4327), .B1(n4277), .B2(n657), .ZN(U57_Z_11)
         );
  OAI22_X2 U883 ( .A1(n719), .A2(n4325), .B1(n4278), .B2(n575), .ZN(U57_Z_109)
         );
  OAI22_X2 U884 ( .A1(n720), .A2(n4325), .B1(n4278), .B2(n576), .ZN(U57_Z_108)
         );
  OAI22_X2 U885 ( .A1(n721), .A2(n4325), .B1(n4278), .B2(n577), .ZN(U57_Z_107)
         );
  OAI22_X2 U886 ( .A1(n722), .A2(n4325), .B1(n4278), .B2(n578), .ZN(U57_Z_106)
         );
  OAI22_X2 U887 ( .A1(n723), .A2(n4325), .B1(n4278), .B2(n579), .ZN(U57_Z_105)
         );
  OAI22_X2 U888 ( .A1(n724), .A2(n4325), .B1(n4278), .B2(n580), .ZN(U57_Z_104)
         );
  OAI22_X2 U889 ( .A1(n725), .A2(n4325), .B1(n4278), .B2(n581), .ZN(U57_Z_103)
         );
  OAI22_X2 U890 ( .A1(n726), .A2(n4325), .B1(n4278), .B2(n582), .ZN(U57_Z_102)
         );
  OAI22_X2 U891 ( .A1(n727), .A2(n4325), .B1(n4278), .B2(n583), .ZN(U57_Z_101)
         );
  OAI22_X2 U892 ( .A1(n728), .A2(n4325), .B1(n4278), .B2(n584), .ZN(U57_Z_100)
         );
  NOR3_X2 U893 ( .A1(n1197), .A2(n1196), .A3(n1192), .ZN(n1198) );
  OAI22_X2 U894 ( .A1(n754), .A2(n4327), .B1(n4277), .B2(n658), .ZN(U57_Z_10)
         );
  OAI22_X2 U895 ( .A1(n763), .A2(n4327), .B1(n4277), .B2(n667), .ZN(U57_Z_1)
         );
  OAI22_X2 U896 ( .A1(n764), .A2(n4327), .B1(n4277), .B2(n668), .ZN(U57_Z_0)
         );
  NAND3_X2 U898 ( .A1(n280), .A2(n1191), .A3(n281), .ZN(n1199) );
  NOR4_X2 U899 ( .A1(n285), .A2(n282), .A3(n283), .A4(n1143), .ZN(n1192) );
  NAND4_X2 U900 ( .A1(n1133), .A2(n1138), .A3(n1143), .A4(n283), .ZN(n1191) );
  NOR4_X2 U901 ( .A1(n282), .A2(n284), .A3(n283), .A4(n1133), .ZN(n1197) );
  NOR4_X2 U903 ( .A1(n285), .A2(n284), .A3(n283), .A4(n1138), .ZN(n1196) );
  NAND2_X2 U908 ( .A1(n1200), .A2(n122), .ZN(U55_Z_1) );
  NAND3_X2 U909 ( .A1(n[3036]), .A2(n125), .A3(n4287), .ZN(n1200) );
  NOR2_X2 U911 ( .A1(n1079), .A2(n123), .ZN(n1127) );
  NOR4_X2 U913 ( .A1(n1206), .A2(n1207), .A3(n1208), .A4(n1209), .ZN(n1205) );
  XOR2_X2 U914 ( .A(n1162), .B(n1178), .Z(n1209) );
  NAND2_X2 U916 ( .A1(n1210), .A2(n124), .ZN(n1162) );
  OAI22_X2 U917 ( .A1(n305), .A2(n4317), .B1(n4320), .B2(n294), .ZN(n1210) );
  XOR2_X2 U918 ( .A(n1158), .B(n1176), .Z(n1208) );
  NAND2_X2 U920 ( .A1(n1211), .A2(n124), .ZN(n1158) );
  OAI22_X2 U921 ( .A1(n303), .A2(n4269), .B1(n4320), .B2(n292), .ZN(n1211) );
  XOR2_X2 U922 ( .A(n1160), .B(n1177), .Z(n1207) );
  NAND2_X2 U924 ( .A1(n1212), .A2(n124), .ZN(n1160) );
  OAI22_X2 U925 ( .A1(n304), .A2(n4317), .B1(n4320), .B2(n293), .ZN(n1212) );
  NAND3_X2 U926 ( .A1(n1213), .A2(n1214), .A3(n1215), .ZN(n1206) );
  XNOR2_X2 U927 ( .A(n1168), .B(n1180), .ZN(n1215) );
  NAND2_X2 U929 ( .A1(n1216), .A2(n124), .ZN(n1168) );
  OAI22_X2 U930 ( .A1(n307), .A2(n4317), .B1(n4320), .B2(n296), .ZN(n1216) );
  XNOR2_X2 U931 ( .A(n1164), .B(n1179), .ZN(n1214) );
  NAND2_X2 U933 ( .A1(n1217), .A2(n124), .ZN(n1164) );
  OAI22_X2 U934 ( .A1(n306), .A2(n4269), .B1(n4320), .B2(n295), .ZN(n1217) );
  XNOR2_X2 U935 ( .A(n1181), .B(n1170), .ZN(n1213) );
  NAND2_X2 U936 ( .A1(n1218), .A2(n124), .ZN(n1170) );
  OAI22_X2 U937 ( .A1(n308), .A2(n4317), .B1(n4320), .B2(n297), .ZN(n1218) );
  NOR3_X2 U939 ( .A1(n1219), .A2(n1220), .A3(n1221), .ZN(n1204) );
  XOR2_X2 U940 ( .A(n1156), .B(n1175), .Z(n1221) );
  NAND2_X2 U942 ( .A1(n1222), .A2(n124), .ZN(n1156) );
  OAI22_X2 U943 ( .A1(n302), .A2(n4317), .B1(n4320), .B2(n291), .ZN(n1222) );
  XOR2_X2 U944 ( .A(n1152), .B(n1174), .Z(n1220) );
  NAND2_X2 U946 ( .A1(n1223), .A2(n124), .ZN(n1152) );
  OAI22_X2 U947 ( .A1(n300), .A2(n4318), .B1(n4320), .B2(n289), .ZN(n1223) );
  XOR2_X2 U948 ( .A(n1153), .B(n1154), .Z(n1219) );
  NAND2_X2 U949 ( .A1(n1224), .A2(n124), .ZN(n1154) );
  OAI22_X2 U950 ( .A1(n301), .A2(n4318), .B1(n4320), .B2(n290), .ZN(n1224) );
  XNOR2_X2 U952 ( .A(n1150), .B(n1148), .ZN(n1203) );
  NAND2_X2 U954 ( .A1(n1225), .A2(n124), .ZN(n1150) );
  OAI22_X2 U955 ( .A1(n299), .A2(n4269), .B1(n4320), .B2(n288), .ZN(n1225) );
  XNOR2_X2 U956 ( .A(n1166), .B(n1165), .ZN(n1202) );
  NAND2_X2 U958 ( .A1(n1226), .A2(n124), .ZN(n1166) );
  OAI22_X2 U960 ( .A1(n298), .A2(n4317), .B1(n4320), .B2(n287), .ZN(n1226) );
  NOR2_X2 U962 ( .A1(n4290), .A2(n772), .ZN(n1171) );
  NOR2_X2 U963 ( .A1(n120), .A2(n4295), .ZN(n1172) );
  NAND2_X2 U965 ( .A1(n[3037]), .A2(n[3036]), .ZN(n778) );
  NAND2_X2 U966 ( .A1(n4287), .A2(n1227), .ZN(n1079) );
  NOR2_X2 U967 ( .A1(n125), .A2(n[3036]), .ZN(n1227) );
  INV_X4 U969 ( .A(n1171), .ZN(n5) );
  INV_X4 U971 ( .A(n1100), .ZN(n7) );
  INV_X4 U972 ( .A(n1099), .ZN(n8) );
  INV_X4 U973 ( .A(n1098), .ZN(n9) );
  INV_X4 U974 ( .A(n1097), .ZN(n10) );
  INV_X4 U975 ( .A(n1096), .ZN(n11) );
  INV_X4 U976 ( .A(n1095), .ZN(n12) );
  INV_X4 U977 ( .A(n1094), .ZN(n13) );
  INV_X4 U978 ( .A(n1093), .ZN(n14) );
  INV_X4 U979 ( .A(n1091), .ZN(n15) );
  INV_X4 U980 ( .A(n1090), .ZN(n16) );
  INV_X4 U981 ( .A(n1089), .ZN(n17) );
  INV_X4 U982 ( .A(n1088), .ZN(n18) );
  INV_X4 U983 ( .A(n1087), .ZN(n19) );
  INV_X4 U984 ( .A(n1086), .ZN(n20) );
  INV_X4 U985 ( .A(n1085), .ZN(n21) );
  INV_X4 U986 ( .A(n1084), .ZN(n22) );
  INV_X4 U987 ( .A(n1017), .ZN(n23) );
  INV_X4 U988 ( .A(n1016), .ZN(n24) );
  INV_X4 U989 ( .A(n1015), .ZN(n25) );
  INV_X4 U990 ( .A(n1014), .ZN(n26) );
  INV_X4 U991 ( .A(n1012), .ZN(n27) );
  INV_X4 U992 ( .A(n1011), .ZN(n28) );
  INV_X4 U993 ( .A(n1010), .ZN(n29) );
  INV_X4 U994 ( .A(n1009), .ZN(n30) );
  INV_X4 U995 ( .A(n1008), .ZN(n31) );
  INV_X4 U996 ( .A(n1007), .ZN(n32) );
  INV_X4 U997 ( .A(n1006), .ZN(n33) );
  INV_X4 U998 ( .A(n1005), .ZN(n34) );
  INV_X4 U999 ( .A(n1004), .ZN(n35) );
  INV_X4 U1000 ( .A(n1003), .ZN(n36) );
  INV_X4 U1001 ( .A(n1001), .ZN(n37) );
  INV_X4 U1002 ( .A(n1000), .ZN(n38) );
  INV_X4 U1003 ( .A(n988), .ZN(n39) );
  INV_X4 U1004 ( .A(n987), .ZN(n40) );
  INV_X4 U1005 ( .A(n986), .ZN(n41) );
  INV_X4 U1006 ( .A(n985), .ZN(n42) );
  INV_X4 U1007 ( .A(n984), .ZN(n43) );
  INV_X4 U1008 ( .A(n983), .ZN(n44) );
  INV_X4 U1009 ( .A(n982), .ZN(n45) );
  INV_X4 U1010 ( .A(n981), .ZN(n46) );
  INV_X4 U1011 ( .A(n978), .ZN(n47) );
  INV_X4 U1012 ( .A(n977), .ZN(n48) );
  INV_X4 U1013 ( .A(n976), .ZN(n49) );
  INV_X4 U1014 ( .A(n975), .ZN(n50) );
  INV_X4 U1015 ( .A(n974), .ZN(n51) );
  INV_X4 U1016 ( .A(n973), .ZN(n52) );
  INV_X4 U1017 ( .A(n972), .ZN(n53) );
  INV_X4 U1018 ( .A(n971), .ZN(n54) );
  INV_X4 U1019 ( .A(n970), .ZN(n55) );
  INV_X4 U1020 ( .A(n969), .ZN(n56) );
  INV_X4 U1021 ( .A(n967), .ZN(n57) );
  INV_X4 U1022 ( .A(n966), .ZN(n58) );
  INV_X4 U1023 ( .A(n965), .ZN(n59) );
  INV_X4 U1024 ( .A(n964), .ZN(n60) );
  INV_X4 U1025 ( .A(n963), .ZN(n61) );
  INV_X4 U1026 ( .A(n962), .ZN(n62) );
  INV_X4 U1027 ( .A(n961), .ZN(n63) );
  INV_X4 U1028 ( .A(n960), .ZN(n64) );
  INV_X4 U1029 ( .A(n959), .ZN(n65) );
  INV_X4 U1030 ( .A(n958), .ZN(n66) );
  INV_X4 U1031 ( .A(n956), .ZN(n67) );
  INV_X4 U1032 ( .A(n955), .ZN(n68) );
  INV_X4 U1033 ( .A(n954), .ZN(n69) );
  INV_X4 U1034 ( .A(n953), .ZN(n70) );
  INV_X4 U1035 ( .A(n952), .ZN(n71) );
  INV_X4 U1036 ( .A(n951), .ZN(n72) );
  INV_X4 U1037 ( .A(n950), .ZN(n73) );
  INV_X4 U1038 ( .A(n949), .ZN(n74) );
  INV_X4 U1039 ( .A(n948), .ZN(n75) );
  INV_X4 U1040 ( .A(n947), .ZN(n76) );
  INV_X4 U1041 ( .A(n945), .ZN(n77) );
  INV_X4 U1042 ( .A(n944), .ZN(n78) );
  INV_X4 U1043 ( .A(n943), .ZN(n79) );
  INV_X4 U1044 ( .A(n942), .ZN(n80) );
  INV_X4 U1045 ( .A(n941), .ZN(n81) );
  INV_X4 U1046 ( .A(n940), .ZN(n82) );
  INV_X4 U1047 ( .A(n939), .ZN(n83) );
  INV_X4 U1048 ( .A(n938), .ZN(n84) );
  INV_X4 U1049 ( .A(n937), .ZN(n85) );
  INV_X4 U1050 ( .A(n934), .ZN(n86) );
  INV_X4 U1051 ( .A(n932), .ZN(n87) );
  INV_X4 U1052 ( .A(n931), .ZN(n88) );
  INV_X4 U1053 ( .A(n930), .ZN(n89) );
  INV_X4 U1054 ( .A(n929), .ZN(n90) );
  INV_X4 U1055 ( .A(n928), .ZN(n91) );
  INV_X4 U1056 ( .A(n927), .ZN(n92) );
  INV_X4 U1057 ( .A(n926), .ZN(n93) );
  INV_X4 U1058 ( .A(n925), .ZN(n94) );
  INV_X4 U1059 ( .A(n924), .ZN(n95) );
  INV_X4 U1060 ( .A(n923), .ZN(n96) );
  INV_X4 U1061 ( .A(n921), .ZN(n97) );
  INV_X4 U1062 ( .A(n920), .ZN(n98) );
  INV_X4 U1063 ( .A(n919), .ZN(n99) );
  INV_X4 U1064 ( .A(n918), .ZN(n100) );
  INV_X4 U1065 ( .A(n917), .ZN(n101) );
  INV_X4 U1066 ( .A(n916), .ZN(n102) );
  INV_X4 U1067 ( .A(n879), .ZN(n103) );
  INV_X4 U1068 ( .A(n878), .ZN(n104) );
  INV_X4 U1069 ( .A(n876), .ZN(n105) );
  INV_X4 U1070 ( .A(n875), .ZN(n106) );
  INV_X4 U1071 ( .A(n874), .ZN(n107) );
  INV_X4 U1072 ( .A(n873), .ZN(n108) );
  INV_X4 U1073 ( .A(n872), .ZN(n109) );
  INV_X4 U1074 ( .A(n871), .ZN(n110) );
  INV_X4 U1075 ( .A(n870), .ZN(n111) );
  INV_X4 U1076 ( .A(n869), .ZN(n112) );
  INV_X4 U1077 ( .A(n868), .ZN(n113) );
  INV_X4 U1078 ( .A(n867), .ZN(n114) );
  INV_X4 U1079 ( .A(n865), .ZN(n115) );
  INV_X4 U1080 ( .A(n864), .ZN(n116) );
  INV_X4 U1081 ( .A(n863), .ZN(n117) );
  INV_X4 U1082 ( .A(n860), .ZN(n118) );
  INV_X4 U1083 ( .A(n773), .ZN(n119) );
  INV_X4 U1084 ( .A(n1079), .ZN(n120) );
  INV_X4 U1085 ( .A(U55_Z_1), .ZN(n121) );
  INV_X4 U1086 ( .A(n1127), .ZN(n122) );
  INV_X4 U1087 ( .A(n992), .ZN(n123) );
  INV_X4 U1089 ( .A(n1077), .ZN(n270) );
  INV_X4 U1090 ( .A(n1121), .ZN(n271) );
  INV_X4 U1091 ( .A(n999), .ZN(n272) );
  INV_X4 U1092 ( .A(n1136), .ZN(n273) );
  INV_X4 U1093 ( .A(n1123), .ZN(n274) );
  INV_X4 U1094 ( .A(n1078), .ZN(n275) );
  INV_X4 U1095 ( .A(n1142), .ZN(n276) );
  INV_X4 U1096 ( .A(n1140), .ZN(n277) );
  INV_X4 U1097 ( .A(n1128), .ZN(n278) );
  INV_X4 U1098 ( .A(n1196), .ZN(n279) );
  INV_X4 U1099 ( .A(n1197), .ZN(n280) );
  INV_X4 U1100 ( .A(n1192), .ZN(n281) );
  INV_X4 U1101 ( .A(n1138), .ZN(n282) );
  INV_X4 U1102 ( .A(n1135), .ZN(n283) );
  INV_X4 U1103 ( .A(n1143), .ZN(n284) );
  INV_X4 U1104 ( .A(n1133), .ZN(n285) );
  INV_X4 U1107 ( .A(cpDoneFlag), .ZN(n445) );
  INV_X4 U1108 ( .A(dpDoneFlag), .ZN(n446) );
  INV_X4 U1109 ( .A(inDiagAddr[10]), .ZN(n447) );
  INV_X4 U1110 ( .A(inDiagAddr[9]), .ZN(n448) );
  INV_X4 U1111 ( .A(inDiagAddr[8]), .ZN(n449) );
  INV_X4 U1112 ( .A(inDiagAddr[7]), .ZN(n450) );
  INV_X4 U1113 ( .A(inDiagAddr[6]), .ZN(n451) );
  INV_X4 U1114 ( .A(inDiagAddr[5]), .ZN(n452) );
  INV_X4 U1115 ( .A(inDiagAddr[4]), .ZN(n453) );
  INV_X4 U1116 ( .A(inDiagAddr[3]), .ZN(n454) );
  INV_X4 U1117 ( .A(inDiagAddr[2]), .ZN(n455) );
  INV_X4 U1118 ( .A(inDiagAddr[1]), .ZN(n456) );
  INV_X4 U1119 ( .A(inDiagAddr[0]), .ZN(n457) );
  INV_X4 U1120 ( .A(inNonDAddr[10]), .ZN(n458) );
  INV_X4 U1121 ( .A(inNonDAddr[9]), .ZN(n459) );
  INV_X4 U1122 ( .A(inNonDAddr[8]), .ZN(n460) );
  INV_X4 U1123 ( .A(inNonDAddr[7]), .ZN(n461) );
  INV_X4 U1124 ( .A(inNonDAddr[6]), .ZN(n462) );
  INV_X4 U1125 ( .A(inNonDAddr[5]), .ZN(n463) );
  INV_X4 U1126 ( .A(inNonDAddr[4]), .ZN(n464) );
  INV_X4 U1127 ( .A(inNonDAddr[3]), .ZN(n465) );
  INV_X4 U1128 ( .A(inNonDAddr[2]), .ZN(n466) );
  INV_X4 U1129 ( .A(inNonDAddr[1]), .ZN(n467) );
  INV_X4 U1130 ( .A(inNonDAddr[0]), .ZN(n468) );
  INV_X4 U1131 ( .A(inDiagOH[3]), .ZN(n469) );
  INV_X4 U1132 ( .A(inDiagOH[2]), .ZN(n470) );
  INV_X4 U1133 ( .A(inDiagOH[1]), .ZN(n471) );
  INV_X4 U1134 ( .A(inDiagOH[0]), .ZN(n472) );
  INV_X4 U1135 ( .A(inNonDiagOH[3]), .ZN(n473) );
  INV_X4 U1136 ( .A(inNonDiagOH[2]), .ZN(n474) );
  INV_X4 U1137 ( .A(inNonDiagOH[1]), .ZN(n475) );
  INV_X4 U1138 ( .A(inNonDiagOH[0]), .ZN(n476) );
  INV_X4 U1139 ( .A(inYreadData2[239]), .ZN(n477) );
  INV_X4 U1140 ( .A(inYreadData2[238]), .ZN(n478) );
  INV_X4 U1141 ( .A(inYreadData2[237]), .ZN(n479) );
  INV_X4 U1142 ( .A(inYreadData2[236]), .ZN(n480) );
  INV_X4 U1143 ( .A(inYreadData2[235]), .ZN(n481) );
  INV_X4 U1144 ( .A(inYreadData2[234]), .ZN(n482) );
  INV_X4 U1145 ( .A(inYreadData2[233]), .ZN(n483) );
  INV_X4 U1146 ( .A(inYreadData2[232]), .ZN(n484) );
  INV_X4 U1147 ( .A(inYreadData2[231]), .ZN(n485) );
  INV_X4 U1148 ( .A(inYreadData2[230]), .ZN(n486) );
  INV_X4 U1149 ( .A(inYreadData2[229]), .ZN(n487) );
  INV_X4 U1150 ( .A(inYreadData2[228]), .ZN(n488) );
  INV_X4 U1151 ( .A(inYreadData2[227]), .ZN(n489) );
  INV_X4 U1152 ( .A(inYreadData2[226]), .ZN(n490) );
  INV_X4 U1153 ( .A(inYreadData2[225]), .ZN(n491) );
  INV_X4 U1154 ( .A(inYreadData2[224]), .ZN(n492) );
  INV_X4 U1155 ( .A(inYreadData2[223]), .ZN(n493) );
  INV_X4 U1156 ( .A(inYreadData2[222]), .ZN(n494) );
  INV_X4 U1157 ( .A(inYreadData2[221]), .ZN(n495) );
  INV_X4 U1158 ( .A(inYreadData2[220]), .ZN(n496) );
  INV_X4 U1159 ( .A(inYreadData2[219]), .ZN(n497) );
  INV_X4 U1160 ( .A(inYreadData2[218]), .ZN(n498) );
  INV_X4 U1161 ( .A(inYreadData2[217]), .ZN(n499) );
  INV_X4 U1162 ( .A(inYreadData2[216]), .ZN(n500) );
  INV_X4 U1163 ( .A(inYreadData2[215]), .ZN(n501) );
  INV_X4 U1164 ( .A(inYreadData2[214]), .ZN(n502) );
  INV_X4 U1165 ( .A(inYreadData2[213]), .ZN(n503) );
  INV_X4 U1166 ( .A(inYreadData2[212]), .ZN(n504) );
  INV_X4 U1167 ( .A(inYreadData2[211]), .ZN(n505) );
  INV_X4 U1168 ( .A(inYreadData2[210]), .ZN(n506) );
  INV_X4 U1169 ( .A(inYreadData2[209]), .ZN(n507) );
  INV_X4 U1170 ( .A(inYreadData2[208]), .ZN(n508) );
  INV_X4 U1171 ( .A(inYreadData2[207]), .ZN(n509) );
  INV_X4 U1172 ( .A(inYreadData2[206]), .ZN(n510) );
  INV_X4 U1173 ( .A(inYreadData2[205]), .ZN(n511) );
  INV_X4 U1174 ( .A(inYreadData2[204]), .ZN(n512) );
  INV_X4 U1175 ( .A(inYreadData2[203]), .ZN(n513) );
  INV_X4 U1176 ( .A(inYreadData2[202]), .ZN(n514) );
  INV_X4 U1177 ( .A(inYreadData2[201]), .ZN(n515) );
  INV_X4 U1178 ( .A(inYreadData2[200]), .ZN(n516) );
  INV_X4 U1179 ( .A(inYreadData2[199]), .ZN(n517) );
  INV_X4 U1180 ( .A(inYreadData2[198]), .ZN(n518) );
  INV_X4 U1181 ( .A(inYreadData2[197]), .ZN(n519) );
  INV_X4 U1182 ( .A(inYreadData2[196]), .ZN(n520) );
  INV_X4 U1183 ( .A(inYreadData2[195]), .ZN(n521) );
  INV_X4 U1184 ( .A(inYreadData2[194]), .ZN(n522) );
  INV_X4 U1185 ( .A(inYreadData2[193]), .ZN(n523) );
  INV_X4 U1186 ( .A(inYreadData2[192]), .ZN(n524) );
  INV_X4 U1187 ( .A(inYreadData2[175]), .ZN(n525) );
  INV_X4 U1188 ( .A(inYreadData2[174]), .ZN(n526) );
  INV_X4 U1189 ( .A(inYreadData2[173]), .ZN(n527) );
  INV_X4 U1190 ( .A(inYreadData2[172]), .ZN(n528) );
  INV_X4 U1191 ( .A(inYreadData2[171]), .ZN(n529) );
  INV_X4 U1192 ( .A(inYreadData2[170]), .ZN(n530) );
  INV_X4 U1193 ( .A(inYreadData2[169]), .ZN(n531) );
  INV_X4 U1194 ( .A(inYreadData2[168]), .ZN(n532) );
  INV_X4 U1195 ( .A(inYreadData2[167]), .ZN(n533) );
  INV_X4 U1196 ( .A(inYreadData2[166]), .ZN(n534) );
  INV_X4 U1197 ( .A(inYreadData2[165]), .ZN(n535) );
  INV_X4 U1198 ( .A(inYreadData2[164]), .ZN(n536) );
  INV_X4 U1199 ( .A(inYreadData2[163]), .ZN(n537) );
  INV_X4 U1200 ( .A(inYreadData2[162]), .ZN(n538) );
  INV_X4 U1201 ( .A(inYreadData2[161]), .ZN(n539) );
  INV_X4 U1202 ( .A(inYreadData2[160]), .ZN(n540) );
  INV_X4 U1203 ( .A(inYreadData2[159]), .ZN(n541) );
  INV_X4 U1204 ( .A(inYreadData2[158]), .ZN(n542) );
  INV_X4 U1205 ( .A(inYreadData2[157]), .ZN(n543) );
  INV_X4 U1206 ( .A(inYreadData2[156]), .ZN(n544) );
  INV_X4 U1207 ( .A(inYreadData2[155]), .ZN(n545) );
  INV_X4 U1208 ( .A(inYreadData2[154]), .ZN(n546) );
  INV_X4 U1209 ( .A(inYreadData2[153]), .ZN(n547) );
  INV_X4 U1210 ( .A(inYreadData2[152]), .ZN(n548) );
  INV_X4 U1211 ( .A(inYreadData2[151]), .ZN(n549) );
  INV_X4 U1212 ( .A(inYreadData2[150]), .ZN(n550) );
  INV_X4 U1213 ( .A(inYreadData2[149]), .ZN(n551) );
  INV_X4 U1214 ( .A(inYreadData2[148]), .ZN(n552) );
  INV_X4 U1215 ( .A(inYreadData2[147]), .ZN(n553) );
  INV_X4 U1216 ( .A(inYreadData2[146]), .ZN(n554) );
  INV_X4 U1217 ( .A(inYreadData2[145]), .ZN(n555) );
  INV_X4 U1218 ( .A(inYreadData2[144]), .ZN(n556) );
  INV_X4 U1219 ( .A(inYreadData2[143]), .ZN(n557) );
  INV_X4 U1220 ( .A(inYreadData2[142]), .ZN(n558) );
  INV_X4 U1221 ( .A(inYreadData2[141]), .ZN(n559) );
  INV_X4 U1222 ( .A(inYreadData2[140]), .ZN(n560) );
  INV_X4 U1223 ( .A(inYreadData2[139]), .ZN(n561) );
  INV_X4 U1224 ( .A(inYreadData2[138]), .ZN(n562) );
  INV_X4 U1225 ( .A(inYreadData2[137]), .ZN(n563) );
  INV_X4 U1226 ( .A(inYreadData2[136]), .ZN(n564) );
  INV_X4 U1227 ( .A(inYreadData2[135]), .ZN(n565) );
  INV_X4 U1228 ( .A(inYreadData2[134]), .ZN(n566) );
  INV_X4 U1229 ( .A(inYreadData2[133]), .ZN(n567) );
  INV_X4 U1230 ( .A(inYreadData2[132]), .ZN(n568) );
  INV_X4 U1231 ( .A(inYreadData2[131]), .ZN(n569) );
  INV_X4 U1232 ( .A(inYreadData2[130]), .ZN(n570) );
  INV_X4 U1233 ( .A(inYreadData2[129]), .ZN(n571) );
  INV_X4 U1234 ( .A(inYreadData2[128]), .ZN(n572) );
  INV_X4 U1235 ( .A(inYreadData2[111]), .ZN(n573) );
  INV_X4 U1236 ( .A(inYreadData2[110]), .ZN(n574) );
  INV_X4 U1237 ( .A(inYreadData2[109]), .ZN(n575) );
  INV_X4 U1238 ( .A(inYreadData2[108]), .ZN(n576) );
  INV_X4 U1239 ( .A(inYreadData2[107]), .ZN(n577) );
  INV_X4 U1240 ( .A(inYreadData2[106]), .ZN(n578) );
  INV_X4 U1241 ( .A(inYreadData2[105]), .ZN(n579) );
  INV_X4 U1242 ( .A(inYreadData2[104]), .ZN(n580) );
  INV_X4 U1243 ( .A(inYreadData2[103]), .ZN(n581) );
  INV_X4 U1244 ( .A(inYreadData2[102]), .ZN(n582) );
  INV_X4 U1245 ( .A(inYreadData2[101]), .ZN(n583) );
  INV_X4 U1246 ( .A(inYreadData2[100]), .ZN(n584) );
  INV_X4 U1247 ( .A(inYreadData2[99]), .ZN(n585) );
  INV_X4 U1248 ( .A(inYreadData2[98]), .ZN(n586) );
  INV_X4 U1249 ( .A(inYreadData2[97]), .ZN(n587) );
  INV_X4 U1250 ( .A(inYreadData2[96]), .ZN(n588) );
  INV_X4 U1251 ( .A(inYreadData2[95]), .ZN(n589) );
  INV_X4 U1252 ( .A(inYreadData2[94]), .ZN(n590) );
  INV_X4 U1253 ( .A(inYreadData2[93]), .ZN(n591) );
  INV_X4 U1254 ( .A(inYreadData2[92]), .ZN(n592) );
  INV_X4 U1255 ( .A(inYreadData2[91]), .ZN(n593) );
  INV_X4 U1256 ( .A(inYreadData2[90]), .ZN(n594) );
  INV_X4 U1257 ( .A(inYreadData2[89]), .ZN(n595) );
  INV_X4 U1258 ( .A(inYreadData2[88]), .ZN(n596) );
  INV_X4 U1259 ( .A(inYreadData2[87]), .ZN(n597) );
  INV_X4 U1260 ( .A(inYreadData2[86]), .ZN(n598) );
  INV_X4 U1261 ( .A(inYreadData2[85]), .ZN(n599) );
  INV_X4 U1262 ( .A(inYreadData2[84]), .ZN(n600) );
  INV_X4 U1263 ( .A(inYreadData2[83]), .ZN(n601) );
  INV_X4 U1264 ( .A(inYreadData2[82]), .ZN(n602) );
  INV_X4 U1265 ( .A(inYreadData2[81]), .ZN(n603) );
  INV_X4 U1266 ( .A(inYreadData2[80]), .ZN(n604) );
  INV_X4 U1267 ( .A(inYreadData2[79]), .ZN(n605) );
  INV_X4 U1268 ( .A(inYreadData2[78]), .ZN(n606) );
  INV_X4 U1269 ( .A(inYreadData2[77]), .ZN(n607) );
  INV_X4 U1270 ( .A(inYreadData2[76]), .ZN(n608) );
  INV_X4 U1271 ( .A(inYreadData2[75]), .ZN(n609) );
  INV_X4 U1272 ( .A(inYreadData2[74]), .ZN(n610) );
  INV_X4 U1273 ( .A(inYreadData2[73]), .ZN(n611) );
  INV_X4 U1274 ( .A(inYreadData2[72]), .ZN(n612) );
  INV_X4 U1275 ( .A(inYreadData2[71]), .ZN(n613) );
  INV_X4 U1276 ( .A(inYreadData2[70]), .ZN(n614) );
  INV_X4 U1277 ( .A(inYreadData2[69]), .ZN(n615) );
  INV_X4 U1278 ( .A(inYreadData2[68]), .ZN(n616) );
  INV_X4 U1279 ( .A(inYreadData2[67]), .ZN(n617) );
  INV_X4 U1280 ( .A(inYreadData2[66]), .ZN(n618) );
  INV_X4 U1281 ( .A(inYreadData2[65]), .ZN(n619) );
  INV_X4 U1282 ( .A(inYreadData2[64]), .ZN(n620) );
  INV_X4 U1283 ( .A(inYreadData2[47]), .ZN(n621) );
  INV_X4 U1284 ( .A(inYreadData2[46]), .ZN(n622) );
  INV_X4 U1285 ( .A(inYreadData2[45]), .ZN(n623) );
  INV_X4 U1286 ( .A(inYreadData2[44]), .ZN(n624) );
  INV_X4 U1287 ( .A(inYreadData2[43]), .ZN(n625) );
  INV_X4 U1288 ( .A(inYreadData2[42]), .ZN(n626) );
  INV_X4 U1289 ( .A(inYreadData2[41]), .ZN(n627) );
  INV_X4 U1290 ( .A(inYreadData2[40]), .ZN(n628) );
  INV_X4 U1291 ( .A(inYreadData2[39]), .ZN(n629) );
  INV_X4 U1292 ( .A(inYreadData2[38]), .ZN(n630) );
  INV_X4 U1293 ( .A(inYreadData2[37]), .ZN(n631) );
  INV_X4 U1294 ( .A(inYreadData2[36]), .ZN(n632) );
  INV_X4 U1295 ( .A(inYreadData2[35]), .ZN(n633) );
  INV_X4 U1296 ( .A(inYreadData2[34]), .ZN(n634) );
  INV_X4 U1297 ( .A(inYreadData2[33]), .ZN(n635) );
  INV_X4 U1298 ( .A(inYreadData2[32]), .ZN(n636) );
  INV_X4 U1299 ( .A(inYreadData2[31]), .ZN(n637) );
  INV_X4 U1300 ( .A(inYreadData2[30]), .ZN(n638) );
  INV_X4 U1301 ( .A(inYreadData2[29]), .ZN(n639) );
  INV_X4 U1302 ( .A(inYreadData2[28]), .ZN(n640) );
  INV_X4 U1303 ( .A(inYreadData2[27]), .ZN(n641) );
  INV_X4 U1304 ( .A(inYreadData2[26]), .ZN(n642) );
  INV_X4 U1305 ( .A(inYreadData2[25]), .ZN(n643) );
  INV_X4 U1306 ( .A(inYreadData2[24]), .ZN(n644) );
  INV_X4 U1307 ( .A(inYreadData2[23]), .ZN(n645) );
  INV_X4 U1308 ( .A(inYreadData2[22]), .ZN(n646) );
  INV_X4 U1309 ( .A(inYreadData2[21]), .ZN(n647) );
  INV_X4 U1310 ( .A(inYreadData2[20]), .ZN(n648) );
  INV_X4 U1311 ( .A(inYreadData2[19]), .ZN(n649) );
  INV_X4 U1312 ( .A(inYreadData2[18]), .ZN(n650) );
  INV_X4 U1313 ( .A(inYreadData2[17]), .ZN(n651) );
  INV_X4 U1314 ( .A(inYreadData2[16]), .ZN(n652) );
  INV_X4 U1315 ( .A(inYreadData2[15]), .ZN(n653) );
  INV_X4 U1316 ( .A(inYreadData2[14]), .ZN(n654) );
  INV_X4 U1317 ( .A(inYreadData2[13]), .ZN(n655) );
  INV_X4 U1318 ( .A(inYreadData2[12]), .ZN(n656) );
  INV_X4 U1319 ( .A(inYreadData2[11]), .ZN(n657) );
  INV_X4 U1320 ( .A(inYreadData2[10]), .ZN(n658) );
  INV_X4 U1321 ( .A(inYreadData2[9]), .ZN(n659) );
  INV_X4 U1322 ( .A(inYreadData2[8]), .ZN(n660) );
  INV_X4 U1323 ( .A(inYreadData2[7]), .ZN(n661) );
  INV_X4 U1324 ( .A(inYreadData2[6]), .ZN(n662) );
  INV_X4 U1325 ( .A(inYreadData2[5]), .ZN(n663) );
  INV_X4 U1326 ( .A(inYreadData2[4]), .ZN(n664) );
  INV_X4 U1327 ( .A(inYreadData2[3]), .ZN(n665) );
  INV_X4 U1328 ( .A(inYreadData2[2]), .ZN(n666) );
  INV_X4 U1329 ( .A(inYreadData2[1]), .ZN(n667) );
  INV_X4 U1330 ( .A(inYreadData2[0]), .ZN(n668) );
  INV_X4 U1331 ( .A(inYComputedVal[47]), .ZN(n669) );
  INV_X4 U1332 ( .A(inYComputedVal[46]), .ZN(n670) );
  INV_X4 U1333 ( .A(inYComputedVal[45]), .ZN(n671) );
  INV_X4 U1334 ( .A(inYComputedVal[44]), .ZN(n672) );
  INV_X4 U1335 ( .A(inYComputedVal[43]), .ZN(n673) );
  INV_X4 U1336 ( .A(inYComputedVal[42]), .ZN(n674) );
  INV_X4 U1337 ( .A(inYComputedVal[41]), .ZN(n675) );
  INV_X4 U1338 ( .A(inYComputedVal[40]), .ZN(n676) );
  INV_X4 U1339 ( .A(inYComputedVal[39]), .ZN(n677) );
  INV_X4 U1340 ( .A(inYComputedVal[38]), .ZN(n678) );
  INV_X4 U1341 ( .A(inYComputedVal[37]), .ZN(n679) );
  INV_X4 U1342 ( .A(inYComputedVal[36]), .ZN(n680) );
  INV_X4 U1343 ( .A(inYComputedVal[35]), .ZN(n681) );
  INV_X4 U1344 ( .A(inYComputedVal[34]), .ZN(n682) );
  INV_X4 U1345 ( .A(inYComputedVal[33]), .ZN(n683) );
  INV_X4 U1346 ( .A(inYComputedVal[32]), .ZN(n684) );
  INV_X4 U1347 ( .A(inYComputedVal[31]), .ZN(n685) );
  INV_X4 U1348 ( .A(inYComputedVal[30]), .ZN(n686) );
  INV_X4 U1349 ( .A(inYComputedVal[29]), .ZN(n687) );
  INV_X4 U1350 ( .A(inYComputedVal[28]), .ZN(n688) );
  INV_X4 U1351 ( .A(inYComputedVal[27]), .ZN(n689) );
  INV_X4 U1352 ( .A(inYComputedVal[26]), .ZN(n690) );
  INV_X4 U1353 ( .A(inYComputedVal[25]), .ZN(n691) );
  INV_X4 U1354 ( .A(inYComputedVal[24]), .ZN(n692) );
  INV_X4 U1355 ( .A(inYComputedVal[23]), .ZN(n693) );
  INV_X4 U1356 ( .A(inYComputedVal[22]), .ZN(n694) );
  INV_X4 U1357 ( .A(inYComputedVal[21]), .ZN(n695) );
  INV_X4 U1358 ( .A(inYComputedVal[20]), .ZN(n696) );
  INV_X4 U1359 ( .A(inYComputedVal[19]), .ZN(n697) );
  INV_X4 U1360 ( .A(inYComputedVal[18]), .ZN(n698) );
  INV_X4 U1361 ( .A(inYComputedVal[17]), .ZN(n699) );
  INV_X4 U1362 ( .A(inYComputedVal[16]), .ZN(n700) );
  INV_X4 U1363 ( .A(inYComputedVal[15]), .ZN(n701) );
  INV_X4 U1364 ( .A(inYComputedVal[14]), .ZN(n702) );
  INV_X4 U1365 ( .A(inYComputedVal[13]), .ZN(n703) );
  INV_X4 U1366 ( .A(inYComputedVal[12]), .ZN(n704) );
  INV_X4 U1367 ( .A(inYComputedVal[11]), .ZN(n705) );
  INV_X4 U1368 ( .A(inYComputedVal[10]), .ZN(n706) );
  INV_X4 U1369 ( .A(inYComputedVal[9]), .ZN(n707) );
  INV_X4 U1370 ( .A(inYComputedVal[8]), .ZN(n708) );
  INV_X4 U1371 ( .A(inYComputedVal[7]), .ZN(n709) );
  INV_X4 U1372 ( .A(inYComputedVal[6]), .ZN(n710) );
  INV_X4 U1373 ( .A(inYComputedVal[5]), .ZN(n711) );
  INV_X4 U1374 ( .A(inYComputedVal[4]), .ZN(n712) );
  INV_X4 U1375 ( .A(inYComputedVal[3]), .ZN(n713) );
  INV_X4 U1376 ( .A(inYComputedVal[2]), .ZN(n714) );
  INV_X4 U1377 ( .A(inYComputedVal[1]), .ZN(n715) );
  INV_X4 U1378 ( .A(inYComputedVal[0]), .ZN(n716) );
  INV_X4 U1379 ( .A(inYchngData[47]), .ZN(n717) );
  INV_X4 U1380 ( .A(inYchngData[46]), .ZN(n718) );
  INV_X4 U1381 ( .A(inYchngData[45]), .ZN(n719) );
  INV_X4 U1382 ( .A(inYchngData[44]), .ZN(n720) );
  INV_X4 U1383 ( .A(inYchngData[43]), .ZN(n721) );
  INV_X4 U1384 ( .A(inYchngData[42]), .ZN(n722) );
  INV_X4 U1385 ( .A(inYchngData[41]), .ZN(n723) );
  INV_X4 U1386 ( .A(inYchngData[40]), .ZN(n724) );
  INV_X4 U1387 ( .A(inYchngData[39]), .ZN(n725) );
  INV_X4 U1388 ( .A(inYchngData[38]), .ZN(n726) );
  INV_X4 U1389 ( .A(inYchngData[37]), .ZN(n727) );
  INV_X4 U1390 ( .A(inYchngData[36]), .ZN(n728) );
  INV_X4 U1391 ( .A(inYchngData[35]), .ZN(n729) );
  INV_X4 U1392 ( .A(inYchngData[34]), .ZN(n730) );
  INV_X4 U1393 ( .A(inYchngData[33]), .ZN(n731) );
  INV_X4 U1394 ( .A(inYchngData[32]), .ZN(n732) );
  INV_X4 U1395 ( .A(inYchngData[31]), .ZN(n733) );
  INV_X4 U1396 ( .A(inYchngData[30]), .ZN(n734) );
  INV_X4 U1397 ( .A(inYchngData[29]), .ZN(n735) );
  INV_X4 U1398 ( .A(inYchngData[28]), .ZN(n736) );
  INV_X4 U1399 ( .A(inYchngData[27]), .ZN(n737) );
  INV_X4 U1400 ( .A(inYchngData[26]), .ZN(n738) );
  INV_X4 U1401 ( .A(inYchngData[25]), .ZN(n739) );
  INV_X4 U1402 ( .A(inYchngData[24]), .ZN(n740) );
  INV_X4 U1403 ( .A(inYchngData[23]), .ZN(n741) );
  INV_X4 U1404 ( .A(inYchngData[22]), .ZN(n742) );
  INV_X4 U1405 ( .A(inYchngData[21]), .ZN(n743) );
  INV_X4 U1406 ( .A(inYchngData[20]), .ZN(n744) );
  INV_X4 U1407 ( .A(inYchngData[19]), .ZN(n745) );
  INV_X4 U1408 ( .A(inYchngData[18]), .ZN(n746) );
  INV_X4 U1409 ( .A(inYchngData[17]), .ZN(n747) );
  INV_X4 U1410 ( .A(inYchngData[16]), .ZN(n748) );
  INV_X4 U1411 ( .A(inYchngData[15]), .ZN(n749) );
  INV_X4 U1412 ( .A(inYchngData[14]), .ZN(n750) );
  INV_X4 U1413 ( .A(inYchngData[13]), .ZN(n751) );
  INV_X4 U1414 ( .A(inYchngData[12]), .ZN(n752) );
  INV_X4 U1415 ( .A(inYchngData[11]), .ZN(n753) );
  INV_X4 U1416 ( .A(inYchngData[10]), .ZN(n754) );
  INV_X4 U1417 ( .A(inYchngData[9]), .ZN(n755) );
  INV_X4 U1418 ( .A(inYchngData[8]), .ZN(n756) );
  INV_X4 U1419 ( .A(inYchngData[7]), .ZN(n757) );
  INV_X4 U1420 ( .A(inYchngData[6]), .ZN(n758) );
  INV_X4 U1421 ( .A(inYchngData[5]), .ZN(n759) );
  INV_X4 U1422 ( .A(inYchngData[4]), .ZN(n760) );
  INV_X4 U1423 ( .A(inYchngData[3]), .ZN(n761) );
  INV_X4 U1424 ( .A(inYchngData[2]), .ZN(n762) );
  INV_X4 U1425 ( .A(inYchngData[1]), .ZN(n763) );
  INV_X4 U1426 ( .A(inYchngData[0]), .ZN(n764) );
  OR3_X1 U1431 ( .A1(n996), .A2(n995), .A3(n999), .ZN(n1104) );
  AND2_X1 U1434 ( .A1(inYreadData2[63]), .A2(n1187), .ZN(U57_Z_63) );
  AND2_X1 U1435 ( .A1(inYreadData2[62]), .A2(n4288), .ZN(U57_Z_62) );
  AND2_X1 U1436 ( .A1(inYreadData2[61]), .A2(n1187), .ZN(U57_Z_61) );
  AND2_X1 U1437 ( .A1(inYreadData2[60]), .A2(n4288), .ZN(U57_Z_60) );
  AND2_X1 U1438 ( .A1(inYreadData2[59]), .A2(n1187), .ZN(U57_Z_59) );
  AND2_X1 U1439 ( .A1(inYreadData2[58]), .A2(n4288), .ZN(U57_Z_58) );
  AND2_X1 U1440 ( .A1(inYreadData2[57]), .A2(n1187), .ZN(U57_Z_57) );
  AND2_X1 U1441 ( .A1(inYreadData2[56]), .A2(n4288), .ZN(U57_Z_56) );
  AND2_X1 U1442 ( .A1(inYreadData2[55]), .A2(n1187), .ZN(U57_Z_55) );
  AND2_X1 U1443 ( .A1(inYreadData2[54]), .A2(n4288), .ZN(U57_Z_54) );
  AND2_X1 U1444 ( .A1(inYreadData2[53]), .A2(n1187), .ZN(U57_Z_53) );
  AND2_X1 U1445 ( .A1(inYreadData2[52]), .A2(n4288), .ZN(U57_Z_52) );
  AND2_X1 U1446 ( .A1(inYreadData2[51]), .A2(n1187), .ZN(U57_Z_51) );
  AND2_X1 U1447 ( .A1(inYreadData2[50]), .A2(n4288), .ZN(U57_Z_50) );
  AND2_X1 U1448 ( .A1(inYreadData2[49]), .A2(n1187), .ZN(U57_Z_49) );
  AND2_X1 U1449 ( .A1(inYreadData2[48]), .A2(n4288), .ZN(U57_Z_48) );
  AND2_X1 U1450 ( .A1(inYreadData2[255]), .A2(n1187), .ZN(U57_Z_255) );
  AND2_X1 U1451 ( .A1(inYreadData2[254]), .A2(n4288), .ZN(U57_Z_254) );
  AND2_X1 U1452 ( .A1(inYreadData2[253]), .A2(n1187), .ZN(U57_Z_253) );
  AND2_X1 U1453 ( .A1(inYreadData2[252]), .A2(n4288), .ZN(U57_Z_252) );
  AND2_X1 U1454 ( .A1(inYreadData2[251]), .A2(n1187), .ZN(U57_Z_251) );
  AND2_X1 U1455 ( .A1(inYreadData2[250]), .A2(n4288), .ZN(U57_Z_250) );
  AND2_X1 U1456 ( .A1(inYreadData2[249]), .A2(n1187), .ZN(U57_Z_249) );
  AND2_X1 U1457 ( .A1(inYreadData2[248]), .A2(n4288), .ZN(U57_Z_248) );
  AND2_X1 U1458 ( .A1(inYreadData2[247]), .A2(n1187), .ZN(U57_Z_247) );
  AND2_X1 U1459 ( .A1(inYreadData2[246]), .A2(n4288), .ZN(U57_Z_246) );
  AND2_X1 U1460 ( .A1(inYreadData2[245]), .A2(n1187), .ZN(U57_Z_245) );
  AND2_X1 U1461 ( .A1(inYreadData2[244]), .A2(n4288), .ZN(U57_Z_244) );
  AND2_X1 U1462 ( .A1(inYreadData2[243]), .A2(n1187), .ZN(U57_Z_243) );
  AND2_X1 U1463 ( .A1(inYreadData2[242]), .A2(n4288), .ZN(U57_Z_242) );
  AND2_X1 U1464 ( .A1(inYreadData2[241]), .A2(n1187), .ZN(U57_Z_241) );
  AND2_X1 U1465 ( .A1(inYreadData2[240]), .A2(n4288), .ZN(U57_Z_240) );
  AND2_X1 U1466 ( .A1(inYreadData2[191]), .A2(n1187), .ZN(U57_Z_191) );
  AND2_X1 U1467 ( .A1(inYreadData2[190]), .A2(n4288), .ZN(U57_Z_190) );
  AND2_X1 U1468 ( .A1(inYreadData2[189]), .A2(n1187), .ZN(U57_Z_189) );
  AND2_X1 U1469 ( .A1(inYreadData2[188]), .A2(n4288), .ZN(U57_Z_188) );
  AND2_X1 U1470 ( .A1(inYreadData2[187]), .A2(n1187), .ZN(U57_Z_187) );
  AND2_X1 U1471 ( .A1(inYreadData2[186]), .A2(n4288), .ZN(U57_Z_186) );
  AND2_X1 U1472 ( .A1(inYreadData2[185]), .A2(n1187), .ZN(U57_Z_185) );
  AND2_X1 U1473 ( .A1(inYreadData2[184]), .A2(n4288), .ZN(U57_Z_184) );
  AND2_X1 U1474 ( .A1(inYreadData2[183]), .A2(n1187), .ZN(U57_Z_183) );
  AND2_X1 U1475 ( .A1(inYreadData2[182]), .A2(n4288), .ZN(U57_Z_182) );
  AND2_X1 U1476 ( .A1(inYreadData2[181]), .A2(n1187), .ZN(U57_Z_181) );
  AND2_X1 U1477 ( .A1(inYreadData2[180]), .A2(n4288), .ZN(U57_Z_180) );
  AND2_X1 U1478 ( .A1(inYreadData2[179]), .A2(n1187), .ZN(U57_Z_179) );
  AND2_X1 U1479 ( .A1(inYreadData2[178]), .A2(n4288), .ZN(U57_Z_178) );
  AND2_X1 U1480 ( .A1(inYreadData2[177]), .A2(n1187), .ZN(U57_Z_177) );
  AND2_X1 U1481 ( .A1(inYreadData2[176]), .A2(n4288), .ZN(U57_Z_176) );
  AND2_X1 U1482 ( .A1(inYreadData2[127]), .A2(n1187), .ZN(U57_Z_127) );
  AND2_X1 U1483 ( .A1(inYreadData2[126]), .A2(n4288), .ZN(U57_Z_126) );
  AND2_X1 U1484 ( .A1(inYreadData2[125]), .A2(n1187), .ZN(U57_Z_125) );
  AND2_X1 U1485 ( .A1(inYreadData2[124]), .A2(n4288), .ZN(U57_Z_124) );
  AND2_X1 U1486 ( .A1(inYreadData2[123]), .A2(n1187), .ZN(U57_Z_123) );
  AND2_X1 U1487 ( .A1(inYreadData2[122]), .A2(n4288), .ZN(U57_Z_122) );
  AND2_X1 U1488 ( .A1(inYreadData2[121]), .A2(n1187), .ZN(U57_Z_121) );
  AND2_X1 U1489 ( .A1(inYreadData2[120]), .A2(n4288), .ZN(U57_Z_120) );
  AND2_X1 U1490 ( .A1(inYreadData2[119]), .A2(n1187), .ZN(U57_Z_119) );
  AND2_X1 U1491 ( .A1(inYreadData2[118]), .A2(n4288), .ZN(U57_Z_118) );
  AND2_X1 U1492 ( .A1(inYreadData2[117]), .A2(n1187), .ZN(U57_Z_117) );
  AND2_X1 U1493 ( .A1(inYreadData2[116]), .A2(n4288), .ZN(U57_Z_116) );
  AND2_X1 U1494 ( .A1(inYreadData2[115]), .A2(n1187), .ZN(U57_Z_115) );
  AND2_X1 U1495 ( .A1(inYreadData2[114]), .A2(n4288), .ZN(U57_Z_114) );
  AND2_X1 U1496 ( .A1(inYreadData2[113]), .A2(n1187), .ZN(U57_Z_113) );
  AND2_X1 U1497 ( .A1(inYreadData2[112]), .A2(n4288), .ZN(U57_Z_112) );
  OR2_X1 U1500 ( .A1(n1161), .A2(n777), .ZN(n1178) );
  OR2_X1 U1501 ( .A1(n1157), .A2(n777), .ZN(n1176) );
  OR2_X1 U1502 ( .A1(n1159), .A2(n777), .ZN(n1177) );
  OR2_X1 U1503 ( .A1(n1167), .A2(n777), .ZN(n1180) );
  OR2_X1 U1504 ( .A1(n1163), .A2(n777), .ZN(n1179) );
  OR2_X1 U1505 ( .A1(n1169), .A2(n777), .ZN(n1181) );
  OR2_X1 U1506 ( .A1(n1155), .A2(n777), .ZN(n1175) );
  OR2_X1 U1507 ( .A1(n1151), .A2(n777), .ZN(n1174) );
  OR2_X1 U1508 ( .A1(n[3036]), .A2(n[3037]), .ZN(n772) );
  DFF_X2 tempNonDiagOH2_reg_3_ ( .D(n1327), .CK(clock), .Q(U35_DATA1_3), .QN(
        n343) );
  DFF_X2 tempNonDiagOH2_reg_2_ ( .D(n1326), .CK(clock), .Q(U35_DATA1_2), .QN(
        n344) );
  DFF_X2 tempNonDiagOH2_reg_1_ ( .D(n1325), .CK(clock), .Q(U35_DATA1_1), .QN(
        n345) );
  DFF_X2 tempNonDiagOH2_reg_0_ ( .D(n1324), .CK(clock), .Q(U35_DATA1_0), .QN(
        n346) );
  DFF_X2 tempDiagOH2_reg_0_ ( .D(n1332), .CK(clock), .Q(U36_DATA1_0), .QN(n338) );
  DFF_X2 tempDiagOH2_reg_3_ ( .D(n1335), .CK(clock), .Q(U36_DATA1_3), .QN(n335) );
  DFF_X2 tempDiagOH2_reg_2_ ( .D(n1334), .CK(clock), .Q(U36_DATA1_2), .QN(n336) );
  DFF_X2 tempDiagOH2_reg_1_ ( .D(n1333), .CK(clock), .Q(U36_DATA1_1), .QN(n337) );
  DFF_X2 tempDiagOH1_reg_3_ ( .D(n1339), .CK(clock), .Q(U36_DATA2_3), .QN(n331) );
  DFF_X2 tempDiagOH1_reg_2_ ( .D(n1338), .CK(clock), .Q(U36_DATA2_2), .QN(n332) );
  DFF_X2 tempNonDiagOH1_reg_3_ ( .D(n1331), .CK(clock), .Q(U35_DATA2_3), .QN(
        n339) );
  DFF_X2 tempNonDiagOH1_reg_2_ ( .D(n1330), .CK(clock), .Q(U35_DATA2_2), .QN(
        n340) );
  DFF_X2 tempNonDiagOH1_reg_1_ ( .D(n1329), .CK(clock), .Q(U35_DATA2_1), .QN(
        n341) );
  DFF_X2 tempNonDiagOH1_reg_0_ ( .D(n1328), .CK(clock), .Q(U35_DATA2_0), .QN(
        n342) );
  DFF_X2 tempNonDiagAddr1_reg_10_ ( .D(n1371), .CK(clock), .Q(U41_DATA2_10), 
        .QN(n309) );
  DFF_X2 tempNonDiagAddr1_reg_9_ ( .D(n1370), .CK(clock), .Q(U41_DATA2_9), 
        .QN(n310) );
  DFF_X2 tempNonDiagAddr1_reg_8_ ( .D(n1369), .CK(clock), .Q(U41_DATA2_8), 
        .QN(n311) );
  DFF_X2 tempNonDiagAddr1_reg_7_ ( .D(n1368), .CK(clock), .Q(U41_DATA2_7), 
        .QN(n312) );
  DFF_X2 tempNonDiagAddr1_reg_6_ ( .D(n1367), .CK(clock), .Q(U41_DATA2_6), 
        .QN(n313) );
  DFF_X2 tempNonDiagAddr1_reg_5_ ( .D(n1366), .CK(clock), .Q(U41_DATA2_5), 
        .QN(n314) );
  DFF_X2 tempNonDiagAddr1_reg_4_ ( .D(n1365), .CK(clock), .Q(U41_DATA2_4), 
        .QN(n315) );
  DFF_X2 tempNonDiagAddr1_reg_3_ ( .D(n1364), .CK(clock), .Q(U41_DATA2_3), 
        .QN(n316) );
  DFF_X2 tempNonDiagAddr1_reg_2_ ( .D(n1363), .CK(clock), .Q(U41_DATA2_2), 
        .QN(n317) );
  DFF_X2 tempNonDiagAddr1_reg_1_ ( .D(n1362), .CK(clock), .Q(U41_DATA2_1), 
        .QN(n318) );
  DFF_X2 tempNonDiagAddr1_reg_0_ ( .D(n1361), .CK(clock), .Q(U41_DATA2_0), 
        .QN(n319) );
  DFF_X2 tempDiagOH1_reg_1_ ( .D(n1337), .CK(clock), .Q(U36_DATA2_1), .QN(n333) );
  DFF_X2 tempDiagOH1_reg_0_ ( .D(n1336), .CK(clock), .Q(U36_DATA2_0), .QN(n334) );
  DFF_X2 tempNonDiagAddr2_reg_0_ ( .D(n1384), .CK(clock), .Q(U41_DATA1_0), 
        .QN(n330) );
  DFF_X2 tempNonDiagAddr2_reg_10_ ( .D(n1349), .CK(clock), .Q(U41_DATA1_10), 
        .QN(n320) );
  DFF_X2 tempNonDiagAddr2_reg_9_ ( .D(n1348), .CK(clock), .Q(U41_DATA1_9), 
        .QN(n321) );
  DFF_X2 tempNonDiagAddr2_reg_8_ ( .D(n1347), .CK(clock), .Q(U41_DATA1_8), 
        .QN(n322) );
  DFF_X2 tempNonDiagAddr2_reg_7_ ( .D(n1346), .CK(clock), .Q(U41_DATA1_7), 
        .QN(n323) );
  DFF_X2 tempNonDiagAddr2_reg_6_ ( .D(n1345), .CK(clock), .Q(U41_DATA1_6), 
        .QN(n324) );
  DFF_X2 tempNonDiagAddr2_reg_5_ ( .D(n1344), .CK(clock), .Q(U41_DATA1_5), 
        .QN(n325) );
  DFF_X2 tempNonDiagAddr2_reg_4_ ( .D(n1343), .CK(clock), .Q(U41_DATA1_4), 
        .QN(n326) );
  DFF_X2 tempNonDiagAddr2_reg_3_ ( .D(n1342), .CK(clock), .Q(U41_DATA1_3), 
        .QN(n327) );
  DFF_X2 tempNonDiagAddr2_reg_2_ ( .D(n1341), .CK(clock), .Q(U41_DATA1_2), 
        .QN(n328) );
  DFF_X2 tempNonDiagAddr2_reg_1_ ( .D(n1340), .CK(clock), .Q(U41_DATA1_1), 
        .QN(n329) );
  DFF_X2 current_state_reg_1_ ( .D(U55_Z_1), .CK(clock), .Q(n[3037]), .QN(n125) );
  DFF_X2 tempDataSecond_reg ( .D(n1383), .CK(clock), .Q(n4279), .QN(n4269) );
  AND2_X4 U161 ( .A1(n120), .A2(n989), .ZN(n4265) );
  AND2_X4 U167 ( .A1(n120), .A2(n997), .ZN(n4268) );
  OR2_X4 U174 ( .A1(n1191), .A2(n122), .ZN(n4271) );
  NAND2_X4 U176 ( .A1(n1127), .A2(n1195), .ZN(n4272) );
  NAND2_X4 U178 ( .A1(n1127), .A2(n1190), .ZN(n4273) );
  AND2_X4 U180 ( .A1(n1127), .A2(n995), .ZN(n805) );
  AND2_X4 U182 ( .A1(n120), .A2(n1074), .ZN(n4274) );
  AND2_X4 U184 ( .A1(n120), .A2(n1129), .ZN(n4275) );
  NAND2_X4 U188 ( .A1(n1127), .A2(n1199), .ZN(n4277) );
  OR2_X4 U190 ( .A1(n122), .A2(n1198), .ZN(n4278) );
  AND2_X4 U192 ( .A1(n4310), .A2(reset), .ZN(n4280) );
  NAND2_X2 U194 ( .A1(n120), .A2(n1101), .ZN(n4281) );
  AND3_X4 U196 ( .A1(n765), .A2(reset), .A3(n775), .ZN(n4282) );
  AND2_X4 U198 ( .A1(n770), .A2(reset), .ZN(n4283) );
  OR2_X4 U200 ( .A1(n1079), .A2(n1080), .ZN(n4284) );
  OR2_X4 U202 ( .A1(n1079), .A2(n1122), .ZN(n4285) );
  OR2_X4 U204 ( .A1(n778), .A2(n4290), .ZN(n4286) );
  AND2_X4 U206 ( .A1(inModuleEnable), .A2(reset), .ZN(n4287) );
  INV_X4 U208 ( .A(n4293), .ZN(n4294) );
  INV_X4 U210 ( .A(n4280), .ZN(n4308) );
  INV_X4 U212 ( .A(n4280), .ZN(n4309) );
  INV_X4 U214 ( .A(n4305), .ZN(n4304) );
  INV_X4 U216 ( .A(n4281), .ZN(n4300) );
  INV_X4 U218 ( .A(n4281), .ZN(n4301) );
  INV_X4 U220 ( .A(n4285), .ZN(n4307) );
  INV_X4 U222 ( .A(n4284), .ZN(n4292) );
  INV_X4 U224 ( .A(n4303), .ZN(n4302) );
  INV_X4 U230 ( .A(n1018), .ZN(n4293) );
  INV_X4 U232 ( .A(n783), .ZN(n4305) );
  INV_X4 U234 ( .A(n4284), .ZN(n4291) );
  INV_X4 U236 ( .A(n4285), .ZN(n4306) );
  INV_X4 U238 ( .A(n4296), .ZN(n4297) );
  INV_X4 U240 ( .A(n802), .ZN(n4303) );
  INV_X4 U242 ( .A(n4296), .ZN(n4299) );
  INV_X4 U244 ( .A(n4295), .ZN(n4298) );
  INV_X4 U246 ( .A(n4282), .ZN(n4312) );
  INV_X4 U248 ( .A(n4282), .ZN(n4313) );
  INV_X4 U250 ( .A(n4316), .ZN(n4314) );
  INV_X4 U251 ( .A(n4316), .ZN(n4315) );
  INV_X4 U252 ( .A(n4283), .ZN(n4310) );
  INV_X4 U253 ( .A(n4283), .ZN(n4311) );
  OAI21_X2 U254 ( .B1(n1102), .B2(n992), .A(n1103), .ZN(n1101) );
  AOI21_X2 U256 ( .B1(n1191), .B2(n1198), .A(n122), .ZN(n4288) );
  AOI21_X2 U257 ( .B1(n1191), .B2(n1198), .A(n122), .ZN(n1187) );
  OAI21_X2 U258 ( .B1(n994), .B2(n1104), .A(n992), .ZN(n1103) );
  INV_X4 U259 ( .A(n4279), .ZN(n4317) );
  AOI22_X2 U260 ( .A1(n1105), .A2(n123), .B1(n992), .B2(n1104), .ZN(n1120) );
  AOI22_X2 U261 ( .A1(n123), .A2(n274), .B1(n992), .B2(n994), .ZN(n1122) );
  AOI22_X2 U262 ( .A1(n993), .A2(n123), .B1(n992), .B2(n996), .ZN(n1080) );
  INV_X4 U264 ( .A(n4320), .ZN(n4318) );
  OAI21_X2 U265 ( .B1(n4290), .B2(n1174), .A(n1173), .ZN(U59_Z_8) );
  OAI21_X2 U266 ( .B1(n4290), .B2(n1175), .A(n1173), .ZN(U59_Z_6) );
  OAI21_X2 U268 ( .B1(n4290), .B2(n1179), .A(n1173), .ZN(U59_Z_2) );
  OAI21_X2 U269 ( .B1(n4290), .B2(n1180), .A(n1173), .ZN(U59_Z_1) );
  OAI21_X2 U270 ( .B1(n4290), .B2(n1177), .A(n1173), .ZN(U59_Z_4) );
  OAI21_X2 U272 ( .B1(n4290), .B2(n1176), .A(n1173), .ZN(U59_Z_5) );
  OAI21_X2 U274 ( .B1(n4290), .B2(n1178), .A(n1173), .ZN(U59_Z_3) );
  OAI21_X2 U276 ( .B1(n4290), .B2(n1181), .A(n1173), .ZN(U59_Z_0) );
  INV_X4 U278 ( .A(n765), .ZN(n4316) );
  NAND4_X2 U280 ( .A1(n1202), .A2(n1203), .A3(n1204), .A4(n1205), .ZN(n992) );
  INV_X4 U282 ( .A(n777), .ZN(n124) );
  INV_X4 U284 ( .A(n4317), .ZN(n4319) );
  NAND2_X2 U286 ( .A1(n4287), .A2(n1182), .ZN(n1173) );
  AOI211_X2 U288 ( .C1(n1142), .C2(n1143), .A(n278), .B(n282), .ZN(n1132) );
  AOI211_X2 U290 ( .C1(n1136), .C2(n1135), .A(n276), .B(n284), .ZN(n1137) );
  AOI211_X2 U292 ( .C1(n1140), .C2(n1133), .A(n273), .B(n283), .ZN(n1141) );
  AOI211_X2 U294 ( .C1(n1128), .C2(n1138), .A(n277), .B(n285), .ZN(n1145) );
  AOI21_X2 U296 ( .B1(n1143), .B2(n1142), .A(n273), .ZN(n1147) );
  AOI21_X2 U298 ( .B1(n1138), .B2(n1128), .A(n276), .ZN(n1146) );
  AOI21_X2 U300 ( .B1(n1135), .B2(n1136), .A(n277), .ZN(n1134) );
  OAI21_X2 U302 ( .B1(n1165), .B2(n4290), .A(n1173), .ZN(U59_Z_10) );
  OAI21_X2 U304 ( .B1(n1148), .B2(n4290), .A(n1173), .ZN(U59_Z_9) );
  OAI21_X2 U306 ( .B1(n1153), .B2(n4290), .A(n1173), .ZN(U59_Z_7) );
  AOI21_X2 U308 ( .B1(n1133), .B2(n1140), .A(n278), .ZN(n1139) );
  INV_X4 U310 ( .A(n4287), .ZN(n4290) );
  INV_X4 U312 ( .A(reset), .ZN(n4321) );
  OAI21_X2 U314 ( .B1(n773), .B2(n776), .A(reset), .ZN(n765) );
  OAI21_X2 U316 ( .B1(n771), .B2(n772), .A(n119), .ZN(n770) );
  AOI222_X1 U318 ( .A1(U6_DATA3_192), .A2(n4295), .B1(n4268), .B2(n859), .C1(
        inYreadData1[192]), .C2(n4265), .ZN(n988) );
  AOI222_X1 U319 ( .A1(U6_DATA3_193), .A2(n4296), .B1(n4268), .B2(n857), .C1(
        inYreadData1[193]), .C2(n4265), .ZN(n987) );
  AOI222_X1 U320 ( .A1(U6_DATA3_194), .A2(n4295), .B1(n4268), .B2(n855), .C1(
        inYreadData1[194]), .C2(n4265), .ZN(n986) );
  AOI222_X1 U321 ( .A1(U6_DATA3_195), .A2(n4295), .B1(n4268), .B2(n853), .C1(
        inYreadData1[195]), .C2(n4265), .ZN(n985) );
  AOI222_X1 U322 ( .A1(U6_DATA3_196), .A2(n4296), .B1(n4268), .B2(n851), .C1(
        inYreadData1[196]), .C2(n4265), .ZN(n984) );
  AOI222_X1 U323 ( .A1(U6_DATA3_197), .A2(n4296), .B1(n4268), .B2(n849), .C1(
        inYreadData1[197]), .C2(n4265), .ZN(n983) );
  AOI222_X1 U324 ( .A1(U6_DATA3_198), .A2(n4295), .B1(n4268), .B2(n846), .C1(
        inYreadData1[198]), .C2(n4265), .ZN(n982) );
  AOI222_X1 U326 ( .A1(U6_DATA3_199), .A2(n4295), .B1(n4268), .B2(n844), .C1(
        inYreadData1[199]), .C2(n4265), .ZN(n981) );
  AOI222_X1 U327 ( .A1(U6_DATA3_200), .A2(n4296), .B1(n4268), .B2(n828), .C1(
        inYreadData1[200]), .C2(n4265), .ZN(n978) );
  AOI222_X1 U328 ( .A1(U6_DATA3_201), .A2(n4295), .B1(n4268), .B2(n806), .C1(
        inYreadData1[201]), .C2(n4265), .ZN(n977) );
  AOI222_X1 U329 ( .A1(U6_DATA3_202), .A2(n4296), .B1(n4268), .B2(n840), .C1(
        inYreadData1[202]), .C2(n4265), .ZN(n976) );
  AOI222_X1 U330 ( .A1(U6_DATA3_203), .A2(n4295), .B1(n4268), .B2(n838), .C1(
        inYreadData1[203]), .C2(n4265), .ZN(n975) );
  AOI22_X2 U331 ( .A1(n4291), .A2(n859), .B1(inYreadData1[128]), .B2(n4323), 
        .ZN(n1073) );
  AOI22_X2 U332 ( .A1(n4291), .A2(n857), .B1(inYreadData1[129]), .B2(n4323), 
        .ZN(n1072) );
  AOI22_X2 U333 ( .A1(n4291), .A2(n855), .B1(inYreadData1[130]), .B2(n4323), 
        .ZN(n1070) );
  AOI22_X2 U334 ( .A1(n4291), .A2(n853), .B1(inYreadData1[131]), .B2(n4323), 
        .ZN(n1069) );
  AOI22_X2 U335 ( .A1(n4291), .A2(n851), .B1(inYreadData1[132]), .B2(n4323), 
        .ZN(n1068) );
  AOI22_X2 U336 ( .A1(n4291), .A2(n849), .B1(inYreadData1[133]), .B2(n4323), 
        .ZN(n1067) );
  AOI22_X2 U338 ( .A1(n4291), .A2(n846), .B1(inYreadData1[134]), .B2(n4323), 
        .ZN(n1066) );
  AOI22_X2 U339 ( .A1(n4291), .A2(n844), .B1(inYreadData1[135]), .B2(n4323), 
        .ZN(n1065) );
  AOI22_X2 U340 ( .A1(n4291), .A2(n828), .B1(inYreadData1[136]), .B2(n4323), 
        .ZN(n1064) );
  AOI22_X2 U341 ( .A1(n4291), .A2(n806), .B1(inYreadData1[137]), .B2(n4323), 
        .ZN(n1063) );
  AOI22_X2 U342 ( .A1(n4291), .A2(n840), .B1(inYreadData1[138]), .B2(n4323), 
        .ZN(n1062) );
  AOI22_X2 U343 ( .A1(n4291), .A2(n838), .B1(inYreadData1[139]), .B2(n4323), 
        .ZN(n1061) );
  AOI22_X2 U344 ( .A1(inYreadData1[26]), .A2(n4275), .B1(n805), .B2(n801), 
        .ZN(n915) );
  AOI22_X2 U345 ( .A1(inYreadData1[27]), .A2(n4275), .B1(n805), .B2(n799), 
        .ZN(n914) );
  AOI22_X2 U346 ( .A1(inYreadData1[28]), .A2(n4275), .B1(n805), .B2(n797), 
        .ZN(n913) );
  AOI22_X2 U347 ( .A1(inYreadData1[29]), .A2(n4275), .B1(n805), .B2(n795), 
        .ZN(n912) );
  AOI22_X2 U348 ( .A1(inYreadData1[30]), .A2(n4275), .B1(n805), .B2(n793), 
        .ZN(n910) );
  AOI22_X2 U350 ( .A1(inYreadData1[31]), .A2(n4275), .B1(n805), .B2(n791), 
        .ZN(n909) );
  AOI22_X2 U351 ( .A1(inYreadData1[1]), .A2(n4275), .B1(n805), .B2(n857), .ZN(
        n1125) );
  AOI22_X2 U352 ( .A1(inYreadData1[10]), .A2(n4275), .B1(n805), .B2(n840), 
        .ZN(n1124) );
  AOI22_X2 U353 ( .A1(n4307), .A2(n840), .B1(inYreadData1[74]), .B2(n4304), 
        .ZN(n839) );
  AOI22_X2 U354 ( .A1(inYreadData1[11]), .A2(n4275), .B1(n805), .B2(n838), 
        .ZN(n1109) );
  AOI22_X2 U355 ( .A1(n4307), .A2(n838), .B1(inYreadData1[75]), .B2(n4304), 
        .ZN(n837) );
  AOI22_X2 U356 ( .A1(inYreadData1[12]), .A2(n4275), .B1(n805), .B2(n836), 
        .ZN(n1092) );
  AOI22_X2 U357 ( .A1(n4307), .A2(n836), .B1(inYreadData1[76]), .B2(n4304), 
        .ZN(n835) );
  AOI22_X2 U358 ( .A1(inYreadData1[13]), .A2(n4275), .B1(n805), .B2(n834), 
        .ZN(n1071) );
  AOI22_X2 U360 ( .A1(inYreadData1[14]), .A2(n4275), .B1(n805), .B2(n832), 
        .ZN(n1060) );
  AOI22_X2 U363 ( .A1(inYreadData1[15]), .A2(n4275), .B1(n805), .B2(n830), 
        .ZN(n1049) );
  AOI22_X2 U364 ( .A1(n4306), .A2(n830), .B1(inYreadData1[79]), .B2(n4304), 
        .ZN(n829) );
  AOI22_X2 U365 ( .A1(inYreadData1[16]), .A2(n4275), .B1(n805), .B2(n826), 
        .ZN(n1038) );
  AOI22_X2 U366 ( .A1(inYreadData1[17]), .A2(n4275), .B1(n805), .B2(n824), 
        .ZN(n1027) );
  AOI22_X2 U367 ( .A1(inYreadData1[18]), .A2(n4275), .B1(n805), .B2(n822), 
        .ZN(n1013) );
  AOI22_X2 U368 ( .A1(inYreadData1[19]), .A2(n4275), .B1(n805), .B2(n820), 
        .ZN(n1002) );
  AOI22_X2 U369 ( .A1(inYreadData1[20]), .A2(n4275), .B1(n805), .B2(n818), 
        .ZN(n979) );
  AOI22_X2 U370 ( .A1(inYreadData1[21]), .A2(n4275), .B1(n805), .B2(n816), 
        .ZN(n968) );
  AOI22_X2 U371 ( .A1(inYreadData1[22]), .A2(n4275), .B1(n805), .B2(n814), 
        .ZN(n957) );
  AOI22_X2 U372 ( .A1(inYreadData1[23]), .A2(n4275), .B1(n805), .B2(n812), 
        .ZN(n946) );
  AOI22_X2 U374 ( .A1(inYreadData1[24]), .A2(n4275), .B1(n805), .B2(n810), 
        .ZN(n933) );
  AOI22_X2 U375 ( .A1(inYreadData1[25]), .A2(n4275), .B1(n805), .B2(n808), 
        .ZN(n922) );
  AOI22_X2 U377 ( .A1(n4307), .A2(n799), .B1(inYreadData1[91]), .B2(n4304), 
        .ZN(n798) );
  AOI22_X2 U379 ( .A1(n4306), .A2(n795), .B1(inYreadData1[93]), .B2(n4304), 
        .ZN(n794) );
  AOI22_X2 U380 ( .A1(n4306), .A2(n793), .B1(inYreadData1[94]), .B2(n783), 
        .ZN(n792) );
  AOI22_X2 U381 ( .A1(n4306), .A2(n791), .B1(inYreadData1[95]), .B2(n783), 
        .ZN(n790) );
  AOI22_X2 U382 ( .A1(inYreadData1[42]), .A2(n4275), .B1(n805), .B2(n891), 
        .ZN(n890) );
  AOI22_X2 U383 ( .A1(inYreadData1[43]), .A2(n4275), .B1(n805), .B2(n889), 
        .ZN(n888) );
  AOI22_X2 U384 ( .A1(inYreadData1[44]), .A2(n4275), .B1(n805), .B2(n887), 
        .ZN(n886) );
  AOI22_X2 U386 ( .A1(inYreadData1[45]), .A2(n4275), .B1(n805), .B2(n885), 
        .ZN(n884) );
  AOI22_X2 U388 ( .A1(inYreadData1[47]), .A2(n4275), .B1(n805), .B2(n881), 
        .ZN(n880) );
  AOI22_X2 U389 ( .A1(inYreadData1[0]), .A2(n4275), .B1(n805), .B2(n859), .ZN(
        n1126) );
  AOI22_X2 U390 ( .A1(inYreadData1[5]), .A2(n4275), .B1(n805), .B2(n849), .ZN(
        n877) );
  AOI22_X2 U391 ( .A1(n4306), .A2(n891), .B1(inYreadData1[106]), .B2(n4304), 
        .ZN(n1113) );
  AOI22_X2 U392 ( .A1(n4306), .A2(n889), .B1(inYreadData1[107]), .B2(n4304), 
        .ZN(n1112) );
  AOI22_X2 U393 ( .A1(n4306), .A2(n887), .B1(inYreadData1[108]), .B2(n4304), 
        .ZN(n1111) );
  AOI22_X2 U394 ( .A1(n4306), .A2(n885), .B1(inYreadData1[109]), .B2(n783), 
        .ZN(n1110) );
  AOI22_X2 U395 ( .A1(n4306), .A2(n883), .B1(inYreadData1[110]), .B2(n783), 
        .ZN(n1108) );
  AOI22_X2 U396 ( .A1(inYreadData1[46]), .A2(n4275), .B1(n805), .B2(n883), 
        .ZN(n882) );
  AOI22_X2 U402 ( .A1(n4306), .A2(n881), .B1(inYreadData1[111]), .B2(n783), 
        .ZN(n1107) );
  AOI22_X2 U403 ( .A1(U36_DATA1_3), .A2(n4279), .B1(n4317), .B2(U36_DATA2_3), 
        .ZN(n1142) );
  AOI21_X2 U405 ( .B1(n125), .B2(n[3036]), .A(n1227), .ZN(n777) );
  AOI22_X2 U406 ( .A1(U41_DATA1_7), .A2(n4319), .B1(n4269), .B2(U41_DATA2_7), 
        .ZN(n1153) );
  AOI22_X2 U407 ( .A1(U41_DATA1_1), .A2(n4319), .B1(n4269), .B2(U41_DATA2_1), 
        .ZN(n1167) );
  AOI22_X2 U408 ( .A1(U41_DATA1_2), .A2(n4319), .B1(n4269), .B2(U41_DATA2_2), 
        .ZN(n1163) );
  AOI22_X2 U409 ( .A1(n4319), .A2(U41_DATA1_0), .B1(n4269), .B2(U41_DATA2_0), 
        .ZN(n1169) );
  AOI22_X2 U410 ( .A1(U41_DATA1_3), .A2(n4319), .B1(n4269), .B2(U41_DATA2_3), 
        .ZN(n1161) );
  AOI22_X2 U411 ( .A1(U41_DATA1_5), .A2(n4319), .B1(n4317), .B2(U41_DATA2_5), 
        .ZN(n1157) );
  AOI22_X2 U412 ( .A1(U41_DATA1_4), .A2(n4319), .B1(n4317), .B2(U41_DATA2_4), 
        .ZN(n1159) );
  AOI22_X2 U413 ( .A1(U41_DATA1_6), .A2(n4319), .B1(n4269), .B2(U41_DATA2_6), 
        .ZN(n1155) );
  AOI22_X2 U414 ( .A1(U41_DATA1_8), .A2(n4319), .B1(n4269), .B2(U41_DATA2_8), 
        .ZN(n1151) );
  AOI22_X2 U415 ( .A1(n4306), .A2(n904), .B1(inYreadData1[100]), .B2(n783), 
        .ZN(n1119) );
  AOI22_X2 U417 ( .A1(n4306), .A2(n902), .B1(inYreadData1[101]), .B2(n783), 
        .ZN(n1118) );
  AOI22_X2 U418 ( .A1(n4306), .A2(n900), .B1(inYreadData1[102]), .B2(n783), 
        .ZN(n1117) );
  AOI22_X2 U419 ( .A1(n4306), .A2(n898), .B1(inYreadData1[103]), .B2(n783), 
        .ZN(n1116) );
  AOI22_X2 U420 ( .A1(n4306), .A2(n895), .B1(inYreadData1[104]), .B2(n783), 
        .ZN(n1115) );
  AOI22_X2 U421 ( .A1(n4306), .A2(n893), .B1(inYreadData1[105]), .B2(n783), 
        .ZN(n1114) );
  AOI22_X2 U423 ( .A1(n4307), .A2(n859), .B1(inYreadData1[64]), .B2(n4304), 
        .ZN(n858) );
  AOI22_X2 U425 ( .A1(n4307), .A2(n857), .B1(inYreadData1[65]), .B2(n4304), 
        .ZN(n856) );
  AOI22_X2 U427 ( .A1(n4307), .A2(n855), .B1(inYreadData1[66]), .B2(n4304), 
        .ZN(n854) );
  AOI22_X2 U429 ( .A1(n4307), .A2(n853), .B1(inYreadData1[67]), .B2(n4304), 
        .ZN(n852) );
  AOI22_X2 U431 ( .A1(n4307), .A2(n851), .B1(inYreadData1[68]), .B2(n4304), 
        .ZN(n850) );
  AOI22_X2 U433 ( .A1(n4307), .A2(n849), .B1(inYreadData1[69]), .B2(n4304), 
        .ZN(n848) );
  AOI22_X2 U435 ( .A1(n4307), .A2(n846), .B1(inYreadData1[70]), .B2(n4304), 
        .ZN(n845) );
  AOI22_X2 U437 ( .A1(n4307), .A2(n844), .B1(inYreadData1[71]), .B2(n4304), 
        .ZN(n843) );
  AOI22_X2 U439 ( .A1(n4307), .A2(n828), .B1(inYreadData1[72]), .B2(n4304), 
        .ZN(n842) );
  AOI22_X2 U441 ( .A1(n4307), .A2(n806), .B1(inYreadData1[73]), .B2(n4304), 
        .ZN(n841) );
  AOI22_X2 U443 ( .A1(n4292), .A2(n836), .B1(inYreadData1[140]), .B2(n4323), 
        .ZN(n1059) );
  AOI22_X2 U445 ( .A1(n4292), .A2(n834), .B1(inYreadData1[141]), .B2(n4323), 
        .ZN(n1058) );
  AOI22_X2 U447 ( .A1(n4292), .A2(n832), .B1(inYreadData1[142]), .B2(n4323), 
        .ZN(n1057) );
  AOI22_X2 U449 ( .A1(n4292), .A2(n830), .B1(inYreadData1[143]), .B2(n4323), 
        .ZN(n1056) );
  AOI22_X2 U452 ( .A1(n4292), .A2(n826), .B1(inYreadData1[144]), .B2(n4323), 
        .ZN(n1055) );
  AOI22_X2 U455 ( .A1(n4306), .A2(n826), .B1(inYreadData1[80]), .B2(n783), 
        .ZN(n825) );
  AOI22_X2 U458 ( .A1(n4292), .A2(n824), .B1(inYreadData1[145]), .B2(n4323), 
        .ZN(n1054) );
  AOI22_X2 U461 ( .A1(n4307), .A2(n824), .B1(inYreadData1[81]), .B2(n4304), 
        .ZN(n823) );
  AOI22_X2 U463 ( .A1(n4292), .A2(n822), .B1(inYreadData1[146]), .B2(n4323), 
        .ZN(n1053) );
  AOI22_X2 U466 ( .A1(n4306), .A2(n822), .B1(inYreadData1[82]), .B2(n4304), 
        .ZN(n821) );
  AOI22_X2 U469 ( .A1(n4292), .A2(n820), .B1(inYreadData1[147]), .B2(n4323), 
        .ZN(n1052) );
  AOI22_X2 U472 ( .A1(n4307), .A2(n820), .B1(inYreadData1[83]), .B2(n783), 
        .ZN(n819) );
  AOI22_X2 U475 ( .A1(n4292), .A2(n818), .B1(inYreadData1[148]), .B2(n4323), 
        .ZN(n1051) );
  AOI22_X2 U478 ( .A1(n4306), .A2(n818), .B1(inYreadData1[84]), .B2(n783), 
        .ZN(n817) );
  AOI22_X2 U481 ( .A1(n4292), .A2(n816), .B1(inYreadData1[149]), .B2(n4323), 
        .ZN(n1050) );
  AOI22_X2 U484 ( .A1(n4307), .A2(n816), .B1(inYreadData1[85]), .B2(n4304), 
        .ZN(n815) );
  AOI22_X2 U487 ( .A1(n4292), .A2(n814), .B1(inYreadData1[150]), .B2(n4323), 
        .ZN(n1048) );
  AOI22_X2 U490 ( .A1(n4307), .A2(n814), .B1(inYreadData1[86]), .B2(n783), 
        .ZN(n813) );
  AOI22_X2 U493 ( .A1(n4292), .A2(n812), .B1(inYreadData1[151]), .B2(n4323), 
        .ZN(n1047) );
  AOI22_X2 U495 ( .A1(n4306), .A2(n812), .B1(inYreadData1[87]), .B2(n4304), 
        .ZN(n811) );
  AOI22_X2 U498 ( .A1(n4292), .A2(n810), .B1(inYreadData1[152]), .B2(n4323), 
        .ZN(n1046) );
  AOI22_X2 U501 ( .A1(n4307), .A2(n810), .B1(inYreadData1[88]), .B2(n783), 
        .ZN(n809) );
  AOI22_X2 U504 ( .A1(n4291), .A2(n808), .B1(inYreadData1[153]), .B2(n4323), 
        .ZN(n1045) );
  AOI22_X2 U507 ( .A1(n4306), .A2(n808), .B1(inYreadData1[89]), .B2(n4304), 
        .ZN(n807) );
  AOI22_X2 U510 ( .A1(n4292), .A2(n801), .B1(inYreadData1[154]), .B2(n4323), 
        .ZN(n1044) );
  AOI22_X2 U513 ( .A1(n4291), .A2(n799), .B1(inYreadData1[155]), .B2(n4323), 
        .ZN(n1043) );
  AOI22_X2 U516 ( .A1(n4292), .A2(n797), .B1(inYreadData1[156]), .B2(n4323), 
        .ZN(n1042) );
  AOI22_X2 U518 ( .A1(n4291), .A2(n795), .B1(inYreadData1[157]), .B2(n4323), 
        .ZN(n1041) );
  AOI22_X2 U520 ( .A1(n4292), .A2(n793), .B1(inYreadData1[158]), .B2(n4323), 
        .ZN(n1040) );
  AOI22_X2 U522 ( .A1(n4291), .A2(n791), .B1(inYreadData1[159]), .B2(n4323), 
        .ZN(n1039) );
  AOI22_X2 U525 ( .A1(n4292), .A2(n789), .B1(inYreadData1[160]), .B2(n4323), 
        .ZN(n1037) );
  AOI22_X2 U527 ( .A1(n4307), .A2(n789), .B1(inYreadData1[96]), .B2(n783), 
        .ZN(n788) );
  AOI22_X2 U529 ( .A1(n4291), .A2(n787), .B1(inYreadData1[161]), .B2(n4323), 
        .ZN(n1036) );
  AOI22_X2 U532 ( .A1(n4306), .A2(n787), .B1(inYreadData1[97]), .B2(n783), 
        .ZN(n786) );
  AOI22_X2 U535 ( .A1(n4292), .A2(n785), .B1(inYreadData1[162]), .B2(n4323), 
        .ZN(n1035) );
  AOI22_X2 U538 ( .A1(n4307), .A2(n785), .B1(inYreadData1[98]), .B2(n783), 
        .ZN(n784) );
  AOI22_X2 U541 ( .A1(n4291), .A2(n782), .B1(inYreadData1[163]), .B2(n4323), 
        .ZN(n1034) );
  AOI22_X2 U544 ( .A1(n4306), .A2(n782), .B1(inYreadData1[99]), .B2(n783), 
        .ZN(n780) );
  AOI22_X2 U547 ( .A1(n4292), .A2(n904), .B1(inYreadData1[164]), .B2(n4323), 
        .ZN(n1033) );
  AOI22_X2 U550 ( .A1(n4291), .A2(n902), .B1(inYreadData1[165]), .B2(n4323), 
        .ZN(n1032) );
  AOI22_X2 U553 ( .A1(n4292), .A2(n900), .B1(inYreadData1[166]), .B2(n4323), 
        .ZN(n1031) );
  AOI22_X2 U556 ( .A1(n4291), .A2(n898), .B1(inYreadData1[167]), .B2(n4323), 
        .ZN(n1030) );
  AOI22_X2 U558 ( .A1(n4291), .A2(n895), .B1(inYreadData1[168]), .B2(n4323), 
        .ZN(n1029) );
  AOI22_X2 U562 ( .A1(n4292), .A2(n893), .B1(inYreadData1[169]), .B2(n4323), 
        .ZN(n1028) );
  AOI22_X2 U563 ( .A1(n4292), .A2(n891), .B1(inYreadData1[170]), .B2(n4323), 
        .ZN(n1026) );
  AOI22_X2 U566 ( .A1(n4291), .A2(n889), .B1(inYreadData1[171]), .B2(n4323), 
        .ZN(n1025) );
  AOI22_X2 U567 ( .A1(n4292), .A2(n887), .B1(inYreadData1[172]), .B2(n4323), 
        .ZN(n1024) );
  AOI22_X2 U568 ( .A1(n4291), .A2(n885), .B1(inYreadData1[173]), .B2(n4323), 
        .ZN(n1023) );
  AOI22_X2 U569 ( .A1(n4291), .A2(n883), .B1(inYreadData1[174]), .B2(n4323), 
        .ZN(n1022) );
  AOI22_X2 U570 ( .A1(n4292), .A2(n881), .B1(inYreadData1[175]), .B2(n4323), 
        .ZN(n1019) );
  AOI22_X2 U571 ( .A1(inYreadData1[2]), .A2(n4275), .B1(n805), .B2(n855), .ZN(
        n980) );
  AOI22_X2 U572 ( .A1(inYreadData1[3]), .A2(n4275), .B1(n805), .B2(n853), .ZN(
        n911) );
  AOI22_X2 U573 ( .A1(inYreadData1[4]), .A2(n4275), .B1(n805), .B2(n851), .ZN(
        n896) );
  AOI22_X2 U575 ( .A1(inYreadData1[6]), .A2(n4275), .B1(n805), .B2(n846), .ZN(
        n866) );
  AOI22_X2 U577 ( .A1(inYreadData1[7]), .A2(n4275), .B1(n805), .B2(n844), .ZN(
        n847) );
  AOI22_X2 U578 ( .A1(inYreadData1[8]), .A2(n4275), .B1(n805), .B2(n828), .ZN(
        n827) );
  AOI22_X2 U579 ( .A1(inYreadData1[9]), .A2(n4275), .B1(n805), .B2(n806), .ZN(
        n803) );
  AOI22_X2 U580 ( .A1(inYreadData1[32]), .A2(n4275), .B1(n805), .B2(n789), 
        .ZN(n908) );
  AOI22_X2 U581 ( .A1(inYreadData1[33]), .A2(n4275), .B1(n805), .B2(n787), 
        .ZN(n907) );
  AOI22_X2 U582 ( .A1(inYreadData1[34]), .A2(n4275), .B1(n805), .B2(n785), 
        .ZN(n906) );
  AOI22_X2 U583 ( .A1(inYreadData1[35]), .A2(n4275), .B1(n805), .B2(n782), 
        .ZN(n905) );
  AOI22_X2 U584 ( .A1(inYreadData1[36]), .A2(n4275), .B1(n805), .B2(n904), 
        .ZN(n903) );
  AOI22_X2 U585 ( .A1(inYreadData1[37]), .A2(n4275), .B1(n805), .B2(n902), 
        .ZN(n901) );
  AOI22_X2 U586 ( .A1(inYreadData1[38]), .A2(n4275), .B1(n805), .B2(n900), 
        .ZN(n899) );
  AOI22_X2 U589 ( .A1(inYreadData1[39]), .A2(n4275), .B1(n805), .B2(n898), 
        .ZN(n897) );
  AOI22_X2 U592 ( .A1(inYreadData1[40]), .A2(n4275), .B1(n805), .B2(n895), 
        .ZN(n894) );
  AOI22_X2 U595 ( .A1(inYreadData1[41]), .A2(n4275), .B1(n805), .B2(n893), 
        .ZN(n892) );
  AOI222_X1 U598 ( .A1(U6_DATA3_204), .A2(n4296), .B1(n4268), .B2(n836), .C1(
        inYreadData1[204]), .C2(n4265), .ZN(n974) );
  AOI222_X1 U601 ( .A1(U6_DATA3_205), .A2(n4296), .B1(n4268), .B2(n834), .C1(
        inYreadData1[205]), .C2(n4265), .ZN(n973) );
  AOI222_X1 U604 ( .A1(U6_DATA3_206), .A2(n4295), .B1(n4268), .B2(n832), .C1(
        inYreadData1[206]), .C2(n4265), .ZN(n972) );
  AOI222_X1 U607 ( .A1(U6_DATA3_207), .A2(n4295), .B1(n4268), .B2(n830), .C1(
        inYreadData1[207]), .C2(n4265), .ZN(n971) );
  AOI222_X1 U610 ( .A1(U6_DATA3_208), .A2(n4296), .B1(n4268), .B2(n826), .C1(
        inYreadData1[208]), .C2(n4265), .ZN(n970) );
  AOI222_X1 U613 ( .A1(U6_DATA3_209), .A2(n4296), .B1(n4268), .B2(n824), .C1(
        inYreadData1[209]), .C2(n4265), .ZN(n969) );
  AOI222_X1 U616 ( .A1(U6_DATA3_210), .A2(n4295), .B1(n4268), .B2(n822), .C1(
        inYreadData1[210]), .C2(n4265), .ZN(n967) );
  AOI222_X1 U619 ( .A1(U6_DATA3_211), .A2(n4295), .B1(n4268), .B2(n820), .C1(
        inYreadData1[211]), .C2(n4265), .ZN(n966) );
  AOI222_X1 U622 ( .A1(U6_DATA3_212), .A2(n4296), .B1(n4268), .B2(n818), .C1(
        inYreadData1[212]), .C2(n4265), .ZN(n965) );
  AOI222_X1 U625 ( .A1(U6_DATA3_213), .A2(n4296), .B1(n4268), .B2(n816), .C1(
        inYreadData1[213]), .C2(n4265), .ZN(n964) );
  AOI222_X1 U627 ( .A1(U6_DATA3_214), .A2(n4295), .B1(n4268), .B2(n814), .C1(
        inYreadData1[214]), .C2(n4265), .ZN(n963) );
  AOI222_X1 U630 ( .A1(U6_DATA3_215), .A2(n4295), .B1(n4268), .B2(n812), .C1(
        inYreadData1[215]), .C2(n4265), .ZN(n962) );
  AOI222_X1 U631 ( .A1(U6_DATA3_216), .A2(n4296), .B1(n4268), .B2(n810), .C1(
        inYreadData1[216]), .C2(n4265), .ZN(n961) );
  AOI222_X1 U632 ( .A1(U6_DATA3_217), .A2(n4295), .B1(n4268), .B2(n808), .C1(
        inYreadData1[217]), .C2(n4265), .ZN(n960) );
  AOI222_X1 U634 ( .A1(U6_DATA3_218), .A2(n4296), .B1(n4268), .B2(n801), .C1(
        inYreadData1[218]), .C2(n4265), .ZN(n959) );
  AOI222_X1 U637 ( .A1(U6_DATA3_219), .A2(n4295), .B1(n4268), .B2(n799), .C1(
        inYreadData1[219]), .C2(n4265), .ZN(n958) );
  AOI222_X1 U640 ( .A1(U6_DATA3_220), .A2(n4296), .B1(n4268), .B2(n797), .C1(
        inYreadData1[220]), .C2(n4265), .ZN(n956) );
  AOI222_X1 U647 ( .A1(U6_DATA3_221), .A2(n4296), .B1(n4268), .B2(n795), .C1(
        inYreadData1[221]), .C2(n4265), .ZN(n955) );
  AOI222_X1 U649 ( .A1(U6_DATA3_222), .A2(n4295), .B1(n4268), .B2(n793), .C1(
        inYreadData1[222]), .C2(n4265), .ZN(n954) );
  AOI222_X1 U651 ( .A1(U6_DATA3_223), .A2(n4296), .B1(n4268), .B2(n791), .C1(
        inYreadData1[223]), .C2(n4265), .ZN(n953) );
  AOI222_X1 U659 ( .A1(U6_DATA3_224), .A2(n4295), .B1(n4268), .B2(n789), .C1(
        inYreadData1[224]), .C2(n4265), .ZN(n952) );
  AOI222_X1 U661 ( .A1(U6_DATA3_225), .A2(n4296), .B1(n4268), .B2(n787), .C1(
        inYreadData1[225]), .C2(n4265), .ZN(n951) );
  AOI222_X1 U662 ( .A1(U6_DATA3_226), .A2(n4295), .B1(n4268), .B2(n785), .C1(
        inYreadData1[226]), .C2(n4265), .ZN(n950) );
  AOI222_X1 U664 ( .A1(U6_DATA3_227), .A2(n4295), .B1(n4268), .B2(n782), .C1(
        inYreadData1[227]), .C2(n4265), .ZN(n949) );
  AOI222_X1 U665 ( .A1(U6_DATA3_228), .A2(n4296), .B1(n4268), .B2(n904), .C1(
        inYreadData1[228]), .C2(n4265), .ZN(n948) );
  AOI222_X1 U666 ( .A1(U6_DATA3_229), .A2(n4296), .B1(n4268), .B2(n902), .C1(
        inYreadData1[229]), .C2(n4265), .ZN(n947) );
  AOI222_X1 U667 ( .A1(U6_DATA3_230), .A2(n4295), .B1(n4268), .B2(n900), .C1(
        inYreadData1[230]), .C2(n4265), .ZN(n945) );
  AOI222_X1 U668 ( .A1(U6_DATA3_231), .A2(n4296), .B1(n4268), .B2(n898), .C1(
        inYreadData1[231]), .C2(n4265), .ZN(n944) );
  AOI222_X1 U669 ( .A1(U6_DATA3_232), .A2(n4295), .B1(n4268), .B2(n895), .C1(
        inYreadData1[232]), .C2(n4265), .ZN(n943) );
  AOI222_X1 U681 ( .A1(U6_DATA3_233), .A2(n4296), .B1(n4268), .B2(n893), .C1(
        inYreadData1[233]), .C2(n4265), .ZN(n942) );
  AOI222_X1 U682 ( .A1(U6_DATA3_234), .A2(n4295), .B1(n4268), .B2(n891), .C1(
        inYreadData1[234]), .C2(n4265), .ZN(n941) );
  AOI222_X1 U683 ( .A1(U6_DATA3_235), .A2(n4295), .B1(n4268), .B2(n889), .C1(
        inYreadData1[235]), .C2(n4265), .ZN(n940) );
  AOI222_X1 U684 ( .A1(U6_DATA3_236), .A2(n4296), .B1(n4268), .B2(n887), .C1(
        inYreadData1[236]), .C2(n4265), .ZN(n939) );
  AOI222_X1 U685 ( .A1(U6_DATA3_237), .A2(n4296), .B1(n4268), .B2(n885), .C1(
        inYreadData1[237]), .C2(n4265), .ZN(n938) );
  AOI222_X1 U686 ( .A1(U6_DATA3_238), .A2(n4295), .B1(n4268), .B2(n883), .C1(
        inYreadData1[238]), .C2(n4265), .ZN(n937) );
  AOI222_X1 U687 ( .A1(U6_DATA3_239), .A2(n4295), .B1(n4268), .B2(n881), .C1(
        inYreadData1[239]), .C2(n4265), .ZN(n934) );
  AOI22_X2 U688 ( .A1(inYreadData1[114]), .A2(n4300), .B1(U6_DATA3_114), .B2(
        n4295), .ZN(n1098) );
  AOI22_X2 U689 ( .A1(inYreadData1[115]), .A2(n4300), .B1(U6_DATA3_115), .B2(
        n4296), .ZN(n1097) );
  AOI22_X2 U690 ( .A1(inYreadData1[50]), .A2(n4300), .B1(U6_DATA3_50), .B2(
        n4296), .ZN(n876) );
  AOI22_X2 U691 ( .A1(inYreadData1[51]), .A2(n4300), .B1(U6_DATA3_51), .B2(
        n4295), .ZN(n875) );
  AOI22_X2 U692 ( .A1(inYreadData1[178]), .A2(n4301), .B1(U6_DATA3_178), .B2(
        n4296), .ZN(n1015) );
  AOI22_X2 U817 ( .A1(inYreadData1[179]), .A2(n4301), .B1(U6_DATA3_179), .B2(
        n4296), .ZN(n1014) );
  AOI22_X2 U819 ( .A1(inYreadData1[240]), .A2(n4301), .B1(U6_DATA3_240), .B2(
        n4295), .ZN(n932) );
  AOI22_X2 U875 ( .A1(inYreadData1[241]), .A2(n4300), .B1(U6_DATA3_241), .B2(
        n4295), .ZN(n931) );
  AOI22_X2 U877 ( .A1(inYreadData1[244]), .A2(n4300), .B1(U6_DATA3_244), .B2(
        n4295), .ZN(n928) );
  AOI22_X2 U879 ( .A1(inYreadData1[245]), .A2(n4301), .B1(U6_DATA3_245), .B2(
        n4296), .ZN(n927) );
  AOI22_X2 U897 ( .A1(inYreadData1[246]), .A2(n4300), .B1(U6_DATA3_246), .B2(
        n4295), .ZN(n926) );
  AOI22_X2 U902 ( .A1(inYreadData1[247]), .A2(n4301), .B1(U6_DATA3_247), .B2(
        n4296), .ZN(n925) );
  AOI22_X2 U904 ( .A1(inYreadData1[242]), .A2(n4301), .B1(U6_DATA3_242), .B2(
        n4296), .ZN(n930) );
  AOI22_X2 U905 ( .A1(inYreadData1[243]), .A2(n4300), .B1(U6_DATA3_243), .B2(
        n4295), .ZN(n929) );
  AOI22_X2 U906 ( .A1(inYreadData1[112]), .A2(n4300), .B1(U6_DATA3_112), .B2(
        n4296), .ZN(n1100) );
  AOI22_X2 U907 ( .A1(inYreadData1[113]), .A2(n4300), .B1(U6_DATA3_113), .B2(
        n4295), .ZN(n1099) );
  AOI22_X2 U910 ( .A1(inYreadData1[116]), .A2(n4300), .B1(U6_DATA3_116), .B2(
        n4295), .ZN(n1096) );
  AOI22_X2 U912 ( .A1(inYreadData1[117]), .A2(n4300), .B1(U6_DATA3_117), .B2(
        n4296), .ZN(n1095) );
  AOI22_X2 U915 ( .A1(inYreadData1[118]), .A2(n4300), .B1(U6_DATA3_118), .B2(
        n4296), .ZN(n1094) );
  AOI22_X2 U919 ( .A1(inYreadData1[119]), .A2(n4300), .B1(U6_DATA3_119), .B2(
        n4295), .ZN(n1093) );
  AOI22_X2 U923 ( .A1(inYreadData1[48]), .A2(n4301), .B1(U6_DATA3_48), .B2(
        n4296), .ZN(n879) );
  AOI22_X2 U928 ( .A1(inYreadData1[49]), .A2(n4300), .B1(U6_DATA3_49), .B2(
        n4295), .ZN(n878) );
  AOI22_X2 U932 ( .A1(inYreadData1[52]), .A2(n4301), .B1(U6_DATA3_52), .B2(
        n4296), .ZN(n874) );
  AOI22_X2 U938 ( .A1(inYreadData1[53]), .A2(n4301), .B1(U6_DATA3_53), .B2(
        n4295), .ZN(n873) );
  AOI22_X2 U941 ( .A1(inYreadData1[54]), .A2(n4300), .B1(U6_DATA3_54), .B2(
        n4296), .ZN(n872) );
  AOI22_X2 U945 ( .A1(inYreadData1[55]), .A2(n4300), .B1(U6_DATA3_55), .B2(
        n4295), .ZN(n871) );
  AOI22_X2 U951 ( .A1(inYreadData1[176]), .A2(n4301), .B1(U6_DATA3_176), .B2(
        n4295), .ZN(n1017) );
  AOI22_X2 U953 ( .A1(inYreadData1[177]), .A2(n4301), .B1(U6_DATA3_177), .B2(
        n4296), .ZN(n1016) );
  AOI22_X2 U957 ( .A1(inYreadData1[180]), .A2(n4301), .B1(U6_DATA3_180), .B2(
        n4296), .ZN(n1012) );
  AOI22_X2 U959 ( .A1(inYreadData1[181]), .A2(n4301), .B1(U6_DATA3_181), .B2(
        n4295), .ZN(n1011) );
  AOI22_X2 U961 ( .A1(inYreadData1[182]), .A2(n4301), .B1(U6_DATA3_182), .B2(
        n4295), .ZN(n1010) );
  AOI22_X2 U964 ( .A1(inYreadData1[183]), .A2(n4301), .B1(U6_DATA3_183), .B2(
        n4296), .ZN(n1009) );
  AOI22_X2 U968 ( .A1(inYreadData1[184]), .A2(n4301), .B1(U6_DATA3_184), .B2(
        n4296), .ZN(n1008) );
  AOI22_X2 U970 ( .A1(inYreadData1[185]), .A2(n4300), .B1(U6_DATA3_185), .B2(
        n4295), .ZN(n1007) );
  AOI22_X2 U1088 ( .A1(inYreadData1[249]), .A2(n4300), .B1(U6_DATA3_249), .B2(
        n4295), .ZN(n923) );
  AOI22_X2 U1105 ( .A1(inYreadData1[248]), .A2(n4301), .B1(U6_DATA3_248), .B2(
        n4296), .ZN(n924) );
  AOI22_X2 U1106 ( .A1(inYreadData1[120]), .A2(n4300), .B1(U6_DATA3_120), .B2(
        n4296), .ZN(n1091) );
  AOI22_X2 U1427 ( .A1(inYreadData1[121]), .A2(n4300), .B1(U6_DATA3_121), .B2(
        n4295), .ZN(n1090) );
  AOI22_X2 U1428 ( .A1(inYreadData1[122]), .A2(n4300), .B1(U6_DATA3_122), .B2(
        n4295), .ZN(n1089) );
  AOI22_X2 U1429 ( .A1(inYreadData1[123]), .A2(n4300), .B1(U6_DATA3_123), .B2(
        n4296), .ZN(n1088) );
  AOI22_X2 U1430 ( .A1(inYreadData1[124]), .A2(n4301), .B1(U6_DATA3_124), .B2(
        n4295), .ZN(n1087) );
  AOI22_X2 U1432 ( .A1(inYreadData1[125]), .A2(n4301), .B1(U6_DATA3_125), .B2(
        n4296), .ZN(n1086) );
  AOI22_X2 U1433 ( .A1(inYreadData1[126]), .A2(n4301), .B1(U6_DATA3_126), .B2(
        n4295), .ZN(n1085) );
  AOI22_X2 U1498 ( .A1(inYreadData1[127]), .A2(n4301), .B1(U6_DATA3_127), .B2(
        n4296), .ZN(n1084) );
  AOI22_X2 U1499 ( .A1(inYreadData1[186]), .A2(n4301), .B1(U6_DATA3_186), .B2(
        n4296), .ZN(n1006) );
  AOI22_X2 U1509 ( .A1(inYreadData1[187]), .A2(n4300), .B1(U6_DATA3_187), .B2(
        n4295), .ZN(n1005) );
  AOI22_X2 U1510 ( .A1(inYreadData1[188]), .A2(n4301), .B1(U6_DATA3_188), .B2(
        n4295), .ZN(n1004) );
  AOI22_X2 U1511 ( .A1(inYreadData1[189]), .A2(n4300), .B1(U6_DATA3_189), .B2(
        n4296), .ZN(n1003) );
  AOI22_X2 U1512 ( .A1(inYreadData1[190]), .A2(n4300), .B1(U6_DATA3_190), .B2(
        n4296), .ZN(n1001) );
  AOI22_X2 U1513 ( .A1(inYreadData1[191]), .A2(n4301), .B1(U6_DATA3_191), .B2(
        n4295), .ZN(n1000) );
  AOI22_X2 U1514 ( .A1(inYreadData1[250]), .A2(n4300), .B1(U6_DATA3_250), .B2(
        n4295), .ZN(n921) );
  AOI22_X2 U1515 ( .A1(inYreadData1[251]), .A2(n4301), .B1(U6_DATA3_251), .B2(
        n4296), .ZN(n920) );
  AOI22_X2 U1516 ( .A1(inYreadData1[252]), .A2(n4300), .B1(U6_DATA3_252), .B2(
        n4295), .ZN(n919) );
  AOI22_X2 U1517 ( .A1(inYreadData1[253]), .A2(n4301), .B1(U6_DATA3_253), .B2(
        n4296), .ZN(n918) );
  AOI22_X2 U1518 ( .A1(inYreadData1[254]), .A2(n4300), .B1(U6_DATA3_254), .B2(
        n4296), .ZN(n917) );
  AOI22_X2 U1519 ( .A1(inYreadData1[255]), .A2(n4301), .B1(U6_DATA3_255), .B2(
        n4295), .ZN(n916) );
  AOI22_X2 U1520 ( .A1(inYreadData1[56]), .A2(n4301), .B1(U6_DATA3_56), .B2(
        n4296), .ZN(n870) );
  AOI22_X2 U1521 ( .A1(inYreadData1[57]), .A2(n4300), .B1(U6_DATA3_57), .B2(
        n4295), .ZN(n869) );
  AOI22_X2 U1522 ( .A1(inYreadData1[58]), .A2(n4301), .B1(U6_DATA3_58), .B2(
        n4295), .ZN(n868) );
  AOI22_X2 U1523 ( .A1(inYreadData1[59]), .A2(n4301), .B1(U6_DATA3_59), .B2(
        n4296), .ZN(n867) );
  AOI22_X2 U1524 ( .A1(inYreadData1[60]), .A2(n4300), .B1(U6_DATA3_60), .B2(
        n4296), .ZN(n865) );
  AOI22_X2 U1525 ( .A1(inYreadData1[61]), .A2(n4300), .B1(U6_DATA3_61), .B2(
        n4295), .ZN(n864) );
  AOI22_X2 U1526 ( .A1(inYreadData1[62]), .A2(n4301), .B1(U6_DATA3_62), .B2(
        n4296), .ZN(n863) );
  AOI22_X2 U1527 ( .A1(inYreadData1[63]), .A2(n4301), .B1(U6_DATA3_63), .B2(
        n4295), .ZN(n860) );
  AOI22_X2 U1528 ( .A1(U35_DATA1_2), .A2(n4319), .B1(n4317), .B2(U35_DATA2_2), 
        .ZN(n1133) );
  AOI22_X2 U1529 ( .A1(U35_DATA1_0), .A2(n4320), .B1(n4317), .B2(U35_DATA2_0), 
        .ZN(n1138) );
  AOI22_X2 U1530 ( .A1(U35_DATA1_3), .A2(n4279), .B1(n4317), .B2(U35_DATA2_3), 
        .ZN(n1143) );
  AOI22_X2 U1531 ( .A1(U35_DATA1_1), .A2(n4279), .B1(n4269), .B2(U35_DATA2_1), 
        .ZN(n1135) );
  AOI22_X2 U1532 ( .A1(U36_DATA1_0), .A2(n4319), .B1(n4269), .B2(U36_DATA2_0), 
        .ZN(n1128) );
  AOI22_X2 U1533 ( .A1(U36_DATA1_1), .A2(n4279), .B1(n4317), .B2(U36_DATA2_1), 
        .ZN(n1136) );
  AOI22_X2 U1534 ( .A1(U36_DATA1_2), .A2(n4319), .B1(n4269), .B2(U36_DATA2_2), 
        .ZN(n1140) );
  AOI22_X2 U1535 ( .A1(U41_DATA1_9), .A2(n4319), .B1(n4269), .B2(U41_DATA2_9), 
        .ZN(n1148) );
  AOI22_X2 U1536 ( .A1(U41_DATA1_10), .A2(n4319), .B1(n4269), .B2(U41_DATA2_10), .ZN(n1165) );
  OAI211_X2 U1537 ( .C1(n4319), .C2(n1172), .A(n1201), .B(n122), .ZN(U55_Z_0)
         );
  OAI21_X2 U1538 ( .B1(n1799), .B2(n4), .A(n1171), .ZN(n1201) );
  NAND3_X2 U1539 ( .A1(n4314), .A2(reset), .A3(n771), .ZN(n4289) );
  INV_X1 U162 ( .A(n4274), .ZN(n4322) );
  INV_X8 U163 ( .A(n4322), .ZN(n4323) );
  INV_X1 U168 ( .A(n4271), .ZN(n4324) );
  INV_X8 U186 ( .A(n4324), .ZN(n4325) );
  INV_X1 U226 ( .A(n4270), .ZN(n4326) );
  INV_X8 U228 ( .A(n4326), .ZN(n4327) );
  NAND2_X2 U263 ( .A1(n1196), .A2(n1127), .ZN(n4270) );
  INV_X1 U297 ( .A(n4267), .ZN(n4328) );
  INV_X8 U299 ( .A(n4328), .ZN(n4329) );
  NAND2_X2 U301 ( .A1(n1192), .A2(n1127), .ZN(n4267) );
  INV_X1 U303 ( .A(n4266), .ZN(n4330) );
  INV_X8 U359 ( .A(n4330), .ZN(n4331) );
  NAND2_X2 U362 ( .A1(n1197), .A2(n1127), .ZN(n4266) );
  OAI221_X1 U376 ( .B1(n717), .B2(n1018), .C1(n4298), .C2(n126), .A(n1019), 
        .ZN(U62_Z_175) );
  OAI221_X1 U378 ( .B1(n718), .B2(n1018), .C1(n4299), .C2(n127), .A(n1022), 
        .ZN(U62_Z_174) );
  OAI221_X1 U422 ( .B1(n719), .B2(n1018), .C1(n4297), .C2(n128), .A(n1023), 
        .ZN(U62_Z_173) );
  OAI221_X1 U424 ( .B1(n720), .B2(n1018), .C1(n4299), .C2(n129), .A(n1024), 
        .ZN(U62_Z_172) );
  AOI22_X1 U426 ( .A1(n4307), .A2(n834), .B1(inYreadData1[77]), .B2(n783), 
        .ZN(n833) );
  AOI22_X1 U428 ( .A1(n4306), .A2(n832), .B1(inYreadData1[78]), .B2(n783), 
        .ZN(n831) );
  AOI22_X1 U1540 ( .A1(n4307), .A2(n801), .B1(inYreadData1[90]), .B2(n783), 
        .ZN(n800) );
  AOI22_X1 U1541 ( .A1(n4307), .A2(n797), .B1(inYreadData1[92]), .B2(n783), 
        .ZN(n796) );
  OAI221_X1 U1542 ( .B1(n729), .B2(n802), .C1(n4297), .C2(n234), .A(n905), 
        .ZN(U62_Z_35) );
  OAI221_X1 U1543 ( .B1(n730), .B2(n802), .C1(n4298), .C2(n235), .A(n906), 
        .ZN(U62_Z_34) );
  OAI221_X1 U1544 ( .B1(n731), .B2(n802), .C1(n4298), .C2(n236), .A(n907), 
        .ZN(U62_Z_33) );
  OAI221_X1 U1545 ( .B1(n732), .B2(n802), .C1(n4286), .C2(n237), .A(n908), 
        .ZN(U62_Z_32) );
  INV_X8 U1546 ( .A(n4286), .ZN(n4295) );
  INV_X8 U1547 ( .A(n4286), .ZN(n4296) );
  INV_X1 U1548 ( .A(n4276), .ZN(n4332) );
  INV_X8 U1549 ( .A(n4332), .ZN(n4333) );
  NAND2_X2 U1550 ( .A1(n1083), .A2(n1106), .ZN(n4276) );
  INV_X8 U1551 ( .A(n4269), .ZN(n4320) );
endmodule


module myDesign ( clock, reset, mydes_chgTxt_row, mydes_chgTxt_col, 
        mydes_chgTxt_real, mydes_chgTxt_img, mydes_ySRAM_rowRead1, 
        mydes_ySRAM_rowRead2, mydes_opYval, mydes_ydataWrite, 
        mydes_op_yReadAddress1, mydes_op_yReadAddress2, mydes_op_yWriteAddress, 
        mydes_op_yWriteEnable, mydes_op_fpIn1, mydes_op_fpIn2, mydes_op_fpMode, 
        mydes_in_fpOut );
  input [15:0] mydes_chgTxt_row;
  input [15:0] mydes_chgTxt_col;
  input [23:0] mydes_chgTxt_real;
  input [23:0] mydes_chgTxt_img;
  input [255:0] mydes_ySRAM_rowRead1;
  input [255:0] mydes_ySRAM_rowRead2;
  output [47:0] mydes_opYval;
  output [255:0] mydes_ydataWrite;
  output [10:0] mydes_op_yReadAddress1;
  output [10:0] mydes_op_yReadAddress2;
  output [10:0] mydes_op_yWriteAddress;
  output [47:0] mydes_op_fpIn1;
  output [47:0] mydes_op_fpIn2;
  input [47:0] mydes_in_fpOut;
  input clock, reset;
  output mydes_op_yWriteEnable, mydes_op_fpMode;
  wire   wire_updateYmoduleEnable, mydes_dataPathDoneFlag, mydes_filtYopDone,
         bWY_op_writeDone, wire_writeYvalEnable, bWY_op_WEbit, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98;
  wire   [10:0] wire_yAddrOut1;
  wire   [10:0] wire_yAddrOut2;
  wire   [10:0] wire_writeDiagAddr;
  wire   [10:0] wire_writeNonDiagAddr;
  wire   [3:0] wire_writeDiagOneHot;
  wire   [3:0] wire_writeNonDiagOneHot;
  wire   [10:0] bWY_op_writeAddress;
  wire   [10:0] bWY_op_readStoreAddr;
  wire   [255:0] bWY_op_writeData;

  updateYcomputation uYc_inst ( .clock(clock), .reset(n97), 
        .computationEnable(wire_updateYmoduleEnable), .uYc_chgTxt_row(
        mydes_chgTxt_row), .uYc_chgTxt_col(mydes_chgTxt_col), 
        .uYc_chgTxt_real(mydes_chgTxt_real), .uYc_chgTxt_img(mydes_chgTxt_img), 
        .uYc_ySRAM_rowRead1(mydes_ySRAM_rowRead1), .uYc_ySRAM_rowRead2(
        mydes_ySRAM_rowRead2), .uYc_yMatAddrOut1(wire_yAddrOut1), 
        .uYc_yMatAddrOut2(wire_yAddrOut2), .uYc_dataPathDoneFlag(
        mydes_dataPathDoneFlag), .uYc_filtYopDone(mydes_filtYopDone), 
        .uYc_opYval(mydes_opYval), .uYc_writeDiagAddr(wire_writeDiagAddr), 
        .uYc_writeNonDiagAddr(wire_writeNonDiagAddr), .uYc_writeDiagOneHot(
        wire_writeDiagOneHot), .uYc_writeNonDiagOneHot(wire_writeNonDiagOneHot), .uYC_op_fpIn1(mydes_op_fpIn1), .uYC_op_fpIn2(mydes_op_fpIn2), 
        .uYC_op_fpMode(mydes_op_fpMode), .uYC_in_fpOut({n96, n94, n92, n90, 
        n88, n86, n84, n82, n80, n78, n76, n74, n72, n70, n68, n66, n64, n62, 
        n60, n58, n56, n54, n52, n50, n48, n46, n44, n42, n40, n38, n36, n34, 
        n32, n30, n28, n26, n24, n22, n20, n18, n16, n14, n12, n10, n8, n6, n4, 
        n2}) );
  roundRobin rR_inst ( .reset(n97), .clock(clock), 
        .in_updateYCtrlPathDoneFlag(mydes_filtYopDone), 
        .in_updateYwriteDoneFlag(bWY_op_writeDone), .op_updateYmoduleEnable(
        wire_updateYmoduleEnable), .op_writeYvalEnable(wire_writeYvalEnable)
         );
  busArbit busArbit_inst ( .reset(n97), .in_yComputeModuleEnable(
        wire_updateYmoduleEnable), .in_yWriteModuleEnable(wire_writeYvalEnable), .in_controlPathReadAddr1(wire_yAddrOut1), .in_controlPathReadAddr2(
        wire_yAddrOut2), .in_controlPathWE(1'b0), .in_controlPathWriteAddr({
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), 
        .in_controlPathWriteData({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .in_writePathReadAddr1(bWY_op_writeAddress), .in_writePathReadAddr2(
        bWY_op_readStoreAddr), .in_writePathWE(bWY_op_WEbit), 
        .in_writePathWriteAddr(bWY_op_writeAddress), .in_writePathWriteData(
        bWY_op_writeData), .op_yReadAddress1(mydes_op_yReadAddress1), 
        .op_yReadAddress2(mydes_op_yReadAddress2), .op_yWriteEnable(
        mydes_op_yWriteEnable), .op_yWriteAddress(mydes_op_yWriteAddress), 
        .op_writeData(mydes_ydataWrite) );
  busWriteY busWriteY_inst ( .clock(clock), .reset(n97), .inModuleEnable(
        wire_writeYvalEnable), .cpDoneFlag(mydes_filtYopDone), .dpDoneFlag(
        mydes_dataPathDoneFlag), .inDiagAddr(wire_writeDiagAddr), .inNonDAddr(
        wire_writeNonDiagAddr), .inDiagOH(wire_writeDiagOneHot), .inNonDiagOH(
        wire_writeNonDiagOneHot), .inYreadData1(mydes_ySRAM_rowRead1), 
        .inYreadData2(mydes_ySRAM_rowRead2), .inYComputedVal(mydes_opYval), 
        .inYchngData({mydes_chgTxt_real, mydes_chgTxt_img}), .op_writeData(
        bWY_op_writeData), .op_writeAddress(bWY_op_writeAddress), 
        .op_readStoreAddr(bWY_op_readStoreAddr), .op_WEbit(bWY_op_WEbit), 
        .op_writeDone(bWY_op_writeDone) );
  INV_X4 U3 ( .A(n98), .ZN(n97) );
  INV_X4 U4 ( .A(reset), .ZN(n98) );
  INV_X4 U5 ( .A(n1), .ZN(n2) );
  INV_X4 U6 ( .A(mydes_in_fpOut[0]), .ZN(n1) );
  INV_X4 U7 ( .A(n3), .ZN(n4) );
  INV_X4 U8 ( .A(mydes_in_fpOut[1]), .ZN(n3) );
  INV_X4 U9 ( .A(n5), .ZN(n6) );
  INV_X4 U10 ( .A(mydes_in_fpOut[2]), .ZN(n5) );
  INV_X4 U11 ( .A(n7), .ZN(n8) );
  INV_X4 U12 ( .A(mydes_in_fpOut[3]), .ZN(n7) );
  INV_X4 U13 ( .A(n9), .ZN(n10) );
  INV_X4 U14 ( .A(mydes_in_fpOut[4]), .ZN(n9) );
  INV_X4 U15 ( .A(n11), .ZN(n12) );
  INV_X4 U16 ( .A(mydes_in_fpOut[5]), .ZN(n11) );
  INV_X4 U17 ( .A(n13), .ZN(n14) );
  INV_X4 U18 ( .A(mydes_in_fpOut[6]), .ZN(n13) );
  INV_X4 U19 ( .A(n15), .ZN(n16) );
  INV_X4 U20 ( .A(mydes_in_fpOut[7]), .ZN(n15) );
  INV_X4 U21 ( .A(n17), .ZN(n18) );
  INV_X4 U22 ( .A(mydes_in_fpOut[8]), .ZN(n17) );
  INV_X4 U23 ( .A(n19), .ZN(n20) );
  INV_X4 U24 ( .A(mydes_in_fpOut[9]), .ZN(n19) );
  INV_X4 U25 ( .A(n21), .ZN(n22) );
  INV_X4 U26 ( .A(mydes_in_fpOut[10]), .ZN(n21) );
  INV_X4 U27 ( .A(n23), .ZN(n24) );
  INV_X4 U28 ( .A(mydes_in_fpOut[11]), .ZN(n23) );
  INV_X4 U29 ( .A(n25), .ZN(n26) );
  INV_X4 U30 ( .A(mydes_in_fpOut[12]), .ZN(n25) );
  INV_X4 U31 ( .A(n27), .ZN(n28) );
  INV_X4 U32 ( .A(mydes_in_fpOut[13]), .ZN(n27) );
  INV_X4 U33 ( .A(n29), .ZN(n30) );
  INV_X4 U34 ( .A(mydes_in_fpOut[14]), .ZN(n29) );
  INV_X4 U35 ( .A(n31), .ZN(n32) );
  INV_X4 U36 ( .A(mydes_in_fpOut[15]), .ZN(n31) );
  INV_X4 U37 ( .A(n33), .ZN(n34) );
  INV_X4 U38 ( .A(mydes_in_fpOut[16]), .ZN(n33) );
  INV_X4 U39 ( .A(n35), .ZN(n36) );
  INV_X4 U40 ( .A(mydes_in_fpOut[17]), .ZN(n35) );
  INV_X4 U41 ( .A(n37), .ZN(n38) );
  INV_X4 U42 ( .A(mydes_in_fpOut[18]), .ZN(n37) );
  INV_X4 U43 ( .A(n39), .ZN(n40) );
  INV_X4 U44 ( .A(mydes_in_fpOut[19]), .ZN(n39) );
  INV_X4 U45 ( .A(n41), .ZN(n42) );
  INV_X4 U46 ( .A(mydes_in_fpOut[20]), .ZN(n41) );
  INV_X4 U47 ( .A(n43), .ZN(n44) );
  INV_X4 U48 ( .A(mydes_in_fpOut[21]), .ZN(n43) );
  INV_X4 U49 ( .A(n45), .ZN(n46) );
  INV_X4 U50 ( .A(mydes_in_fpOut[22]), .ZN(n45) );
  INV_X4 U51 ( .A(n47), .ZN(n48) );
  INV_X4 U52 ( .A(mydes_in_fpOut[23]), .ZN(n47) );
  INV_X4 U53 ( .A(n49), .ZN(n50) );
  INV_X4 U54 ( .A(mydes_in_fpOut[24]), .ZN(n49) );
  INV_X4 U55 ( .A(n51), .ZN(n52) );
  INV_X4 U56 ( .A(mydes_in_fpOut[25]), .ZN(n51) );
  INV_X4 U57 ( .A(n53), .ZN(n54) );
  INV_X4 U58 ( .A(mydes_in_fpOut[26]), .ZN(n53) );
  INV_X4 U59 ( .A(n55), .ZN(n56) );
  INV_X4 U60 ( .A(mydes_in_fpOut[27]), .ZN(n55) );
  INV_X4 U61 ( .A(n57), .ZN(n58) );
  INV_X4 U62 ( .A(mydes_in_fpOut[28]), .ZN(n57) );
  INV_X4 U63 ( .A(n59), .ZN(n60) );
  INV_X4 U64 ( .A(mydes_in_fpOut[29]), .ZN(n59) );
  INV_X4 U65 ( .A(n61), .ZN(n62) );
  INV_X4 U66 ( .A(mydes_in_fpOut[30]), .ZN(n61) );
  INV_X4 U67 ( .A(n63), .ZN(n64) );
  INV_X4 U68 ( .A(mydes_in_fpOut[31]), .ZN(n63) );
  INV_X4 U69 ( .A(n65), .ZN(n66) );
  INV_X4 U70 ( .A(mydes_in_fpOut[32]), .ZN(n65) );
  INV_X4 U71 ( .A(n67), .ZN(n68) );
  INV_X4 U72 ( .A(mydes_in_fpOut[33]), .ZN(n67) );
  INV_X4 U73 ( .A(n69), .ZN(n70) );
  INV_X4 U74 ( .A(mydes_in_fpOut[34]), .ZN(n69) );
  INV_X4 U75 ( .A(n71), .ZN(n72) );
  INV_X4 U76 ( .A(mydes_in_fpOut[35]), .ZN(n71) );
  INV_X4 U77 ( .A(n73), .ZN(n74) );
  INV_X4 U78 ( .A(mydes_in_fpOut[36]), .ZN(n73) );
  INV_X4 U79 ( .A(n75), .ZN(n76) );
  INV_X4 U80 ( .A(mydes_in_fpOut[37]), .ZN(n75) );
  INV_X4 U81 ( .A(n77), .ZN(n78) );
  INV_X4 U82 ( .A(mydes_in_fpOut[38]), .ZN(n77) );
  INV_X4 U83 ( .A(n79), .ZN(n80) );
  INV_X4 U84 ( .A(mydes_in_fpOut[39]), .ZN(n79) );
  INV_X4 U85 ( .A(n81), .ZN(n82) );
  INV_X4 U86 ( .A(mydes_in_fpOut[40]), .ZN(n81) );
  INV_X4 U87 ( .A(n83), .ZN(n84) );
  INV_X4 U88 ( .A(mydes_in_fpOut[41]), .ZN(n83) );
  INV_X4 U89 ( .A(n85), .ZN(n86) );
  INV_X4 U90 ( .A(mydes_in_fpOut[42]), .ZN(n85) );
  INV_X4 U91 ( .A(n87), .ZN(n88) );
  INV_X4 U92 ( .A(mydes_in_fpOut[43]), .ZN(n87) );
  INV_X4 U93 ( .A(n89), .ZN(n90) );
  INV_X4 U94 ( .A(mydes_in_fpOut[44]), .ZN(n89) );
  INV_X4 U95 ( .A(n91), .ZN(n92) );
  INV_X4 U96 ( .A(mydes_in_fpOut[45]), .ZN(n91) );
  INV_X4 U97 ( .A(n93), .ZN(n94) );
  INV_X4 U98 ( .A(mydes_in_fpOut[46]), .ZN(n93) );
  INV_X4 U99 ( .A(n95), .ZN(n96) );
  INV_X4 U100 ( .A(mydes_in_fpOut[47]), .ZN(n95) );
endmodule

