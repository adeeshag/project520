/************************************************************
 *
 * This module is the datapath for the change in Y matrix
 * update. 
 * "Compute_EN" signal so that the Y Computation module does
 * not pull out anymore data. It should sit idle till the next
 * read from change.txt, i.e a computation/ all the iters 
 * should be done.
 *
 * Inputs: 1. Two Y values from the control path. Second value
 *            might be 0 the second read.
 *         2. Execute Enable - module doesn't compute when 0
 *         3. clock,rst
 *    
 * Output: 1. Output of Computation. 
 *            -> this value is not valid if "DoneFlag" is 0
 *         2. DoneFlag - indicates that Computation is done
 *
 * **********************************************************/

module updateY_calc(clock,reset, executeEnableBit,
                     yInVal1, yInVal2, 
                     op_yWriteVal, op_DoneFlag, op_ExDoneFlag
                    );
/* Inputs and Outputs */

input          clock,reset,executeEnableBit;
input [47:0]   yInVal1,yInVal2;

output [47:0]  op_yWriteVal;
output         op_DoneFlag,op_ExDoneFlag;


/* Wires and Regs */
wire        wire_DoneFlag_CmplxMod;

reg [47:0]  op_yWriteVal;
reg         op_DoneFlag,op_ExDoneFlag;

   //Stored in Registers
reg [47:0]  temp_yComputedVal;
reg         temp_nextMode;

   //Wires
reg [47:0] reg_addsubOut;
reg [47:0] reg_addsub_in1,reg_addsub_in2;
 

/* Main Circuit Logic */
always@(posedge clock)
begin
   if(~(reset&executeEnableBit)) // Reset or Enable are 0
   begin
      op_yWriteVal      <= 48'b0;
      op_DoneFlag       <= 1'b0;
      temp_nextMode     <= 1'b1; // always start with subtract first

      temp_yComputedVal <= 48'b0;
      op_ExDoneFlag     <=  1'b0;
      
   end//if-reset
   else
   begin
      if(wire_DoneFlag_CmplxMod) 
      begin
         if(temp_nextMode)
         begin
            op_ExDoneFlag  <= 1'b1;
            temp_nextMode  <= 1'b0; // set to adder next
            op_DoneFlag    <= 1'b0;
            op_yWriteVal   <= 48'b0;
         end
         else // temp_nextMode==0
         begin
            op_yWriteVal   <= reg_addsubOut;
            temp_nextMode  <= 1'b1; // Reset to subtractor next
            op_ExDoneFlag  <= 1'b1;
            op_DoneFlag    <= 1'b1;
         end // temp_nextMode

      end//---if wire_DoneFlag_CmplxMod is high
      else
      begin
         op_yWriteVal   <= 48'b0;
         op_DoneFlag    <= 1'b0;
         op_ExDoneFlag  <= 1'b0;
         // temp_nextMode should retain it's previous value
      end// else wire_DoneFlag_CmplxMod

      temp_yComputedVal <= reg_addsubOut;

   end//-- else-reset

end//posedge clk

      //Deciding inputs and mode to addsub module
always@(*)
begin
   reg_addsub_in1     = yInVal1;

   if(temp_nextMode)
   begin
      reg_addsub_in2  = yInVal2;
   end
   else
   begin
      reg_addsub_in2  = temp_yComputedVal;
   end


end// always@(*)


/* Modules */

addsub_cplx u1 (.clock(clock),.reset(reset),.in1(reg_addsub_in1),.in2(reg_addsub_in2),.mode(temp_nextMode),
                  .op(reg_addsubOut),.done_flag(wire_DoneFlag_CmplxMod),.enable(executeEnableBit)
               );


endmodule




